`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2024 Talha Mahboob
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
///////////////////////////////////////////////////////////////////////////////


//This is the Top Level module for 32-bit Wallace Multiplier
//In this module first we find all the partial products of incoming bits
//Then we add our partial product using Half Adders and Full Adders
//After the Addition of Partial Product we will assign the addition result to our 64-bit Final product

module Wallace_Multiplier_32Bit (
  input  logic [32-1:0] Input1       ,
  input  logic [32-1:0] Input2       ,
  output logic [64-1:0] Final_Product
);

//partial product in the form of array 32x32
  logic [31:0] Partial_Product[31:0];
//Sum and carries generated inter between
  logic [1116:0] Sum      ;
  logic [1116:0] Carry_out;

  genvar i, j;
  generate
    for (i = 0; i < 32; i = i + 1) begin : gen_partial_products
      for (j = 0; j < 32; j = j + 1) begin : gen_bits
        assign Partial_Product[i][j] = Input1[i] & Input2[j];
      end
    end
  endgenerate


//Instantiating Full Adders and Half Adders
//In order to add our partial products
  HalfAdder HA1 (Partial_Product[0][1],Partial_Product[1][0],Sum[0],Carry_out[0]);
  FullAdder FA2 (Partial_Product[0][2],Partial_Product[1][1],Partial_Product[2][0],Sum[1],Carry_out[1]);
  FullAdder FA3 (Partial_Product[0][3],Partial_Product[1][2],Partial_Product[2][1],Sum[2],Carry_out[2]);
  FullAdder FA4 (Partial_Product[0][4],Partial_Product[1][3],Partial_Product[2][2],Sum[3],Carry_out[3]);
  HalfAdder HA5 (Partial_Product[3][1],Partial_Product[4][0],Sum[4],Carry_out[4]);
  FullAdder FA6 (Partial_Product[0][5],Partial_Product[1][4],Partial_Product[2][3],Sum[5],Carry_out[5]);
  FullAdder FA7 (Partial_Product[3][2],Partial_Product[4][1],Partial_Product[5][0],Sum[6],Carry_out[6]);
  FullAdder FA8 (Partial_Product[0][6],Partial_Product[1][5],Partial_Product[2][4],Sum[7],Carry_out[7]);
  FullAdder FA9 (Partial_Product[3][3],Partial_Product[4][2],Partial_Product[5][1],Sum[8],Carry_out[8]);
  FullAdder FA10 (Partial_Product[0][7],Partial_Product[1][6],Partial_Product[2][5],Sum[9],Carry_out[9]);
  FullAdder FA11 (Partial_Product[3][4],Partial_Product[4][3],Partial_Product[5][2],Sum[10],Carry_out[10]);
  HalfAdder HA12 (Partial_Product[6][1],Partial_Product[7][0],Sum[11],Carry_out[11]);
  FullAdder FA13 (Partial_Product[0][8],Partial_Product[1][7],Partial_Product[2][6],Sum[12],Carry_out[12]);
  FullAdder FA14 (Partial_Product[3][5],Partial_Product[4][4],Partial_Product[5][3],Sum[13],Carry_out[13]);
  FullAdder FA15 (Partial_Product[6][2],Partial_Product[7][1],Partial_Product[8][0],Sum[14],Carry_out[14]);
  FullAdder FA16 (Partial_Product[0][9],Partial_Product[1][8],Partial_Product[2][7],Sum[15],Carry_out[15]);
  FullAdder FA17 (Partial_Product[3][6],Partial_Product[4][5],Partial_Product[5][4],Sum[16],Carry_out[16]);
  FullAdder FA18 (Partial_Product[6][3],Partial_Product[7][2],Partial_Product[8][1],Sum[17],Carry_out[17]);
  FullAdder FA19 (Partial_Product[0][10],Partial_Product[1][9],Partial_Product[2][8],Sum[18],Carry_out[18]);
  FullAdder FA20 (Partial_Product[3][7],Partial_Product[4][6],Partial_Product[5][5],Sum[19],Carry_out[19]);
  FullAdder FA21 (Partial_Product[6][4],Partial_Product[7][3],Partial_Product[8][2],Sum[20],Carry_out[20]);
  HalfAdder HA22 (Partial_Product[9][1],Partial_Product[10][0],Sum[21],Carry_out[21]);
  FullAdder FA23 (Partial_Product[0][11],Partial_Product[1][10],Partial_Product[2][9],Sum[22],Carry_out[22]);
  FullAdder FA24 (Partial_Product[3][8],Partial_Product[4][7],Partial_Product[5][6],Sum[23],Carry_out[23]);
  FullAdder FA25 (Partial_Product[6][5],Partial_Product[7][4],Partial_Product[8][3],Sum[24],Carry_out[24]);
  FullAdder FA26 (Partial_Product[9][2],Partial_Product[10][1],Partial_Product[11][0],Sum[25],Carry_out[25]);
  FullAdder FA27 (Partial_Product[0][12],Partial_Product[1][11],Partial_Product[2][10],Sum[26],Carry_out[26]);
  FullAdder FA28 (Partial_Product[3][9],Partial_Product[4][8],Partial_Product[5][7],Sum[27],Carry_out[27]);
  FullAdder FA29 (Partial_Product[6][6],Partial_Product[7][5],Partial_Product[8][4],Sum[28],Carry_out[28]);
  FullAdder FA30 (Partial_Product[9][3],Partial_Product[10][2],Partial_Product[11][1],Sum[29],Carry_out[29]);
  FullAdder FA31 (Partial_Product[0][13],Partial_Product[1][12],Partial_Product[2][11],Sum[30],Carry_out[30]);
  FullAdder FA32 (Partial_Product[3][10],Partial_Product[4][9],Partial_Product[5][8],Sum[31],Carry_out[31]);
  FullAdder FA33 (Partial_Product[6][7],Partial_Product[7][6],Partial_Product[8][5],Sum[32],Carry_out[32]);
  FullAdder FA34 (Partial_Product[9][4],Partial_Product[10][3],Partial_Product[11][2],Sum[33],Carry_out[33]);
  HalfAdder HA35 (Partial_Product[12][1],Partial_Product[13][0],Sum[34],Carry_out[34]);
  FullAdder FA36 (Partial_Product[0][14],Partial_Product[1][13],Partial_Product[2][12],Sum[35],Carry_out[35]);
  FullAdder FA37 (Partial_Product[3][11],Partial_Product[4][10],Partial_Product[5][9],Sum[36],Carry_out[36]);
  FullAdder FA38 (Partial_Product[6][8],Partial_Product[7][7],Partial_Product[8][6],Sum[37],Carry_out[37]);
  FullAdder FA39 (Partial_Product[9][5],Partial_Product[10][4],Partial_Product[11][3],Sum[38],Carry_out[38]);
  FullAdder FA40 (Partial_Product[12][2],Partial_Product[13][1],Partial_Product[14][0],Sum[39],Carry_out[39]);
  FullAdder FA41 (Partial_Product[0][15],Partial_Product[1][14],Partial_Product[2][13],Sum[40],Carry_out[40]);
  FullAdder FA42 (Partial_Product[3][12],Partial_Product[4][11],Partial_Product[5][10],Sum[41],Carry_out[41]);
  FullAdder FA43 (Partial_Product[6][9],Partial_Product[7][8],Partial_Product[8][7],Sum[42],Carry_out[42]);
  FullAdder FA44 (Partial_Product[9][6],Partial_Product[10][5],Partial_Product[11][4],Sum[43],Carry_out[43]);
  FullAdder FA45 (Partial_Product[12][3],Partial_Product[13][2],Partial_Product[14][1],Sum[44],Carry_out[44]);
  FullAdder FA46 (Partial_Product[0][16],Partial_Product[1][15],Partial_Product[2][14],Sum[45],Carry_out[45]);
  FullAdder FA47 (Partial_Product[3][13],Partial_Product[4][12],Partial_Product[5][11],Sum[46],Carry_out[46]);
  FullAdder FA48 (Partial_Product[6][10],Partial_Product[7][9],Partial_Product[8][8],Sum[47],Carry_out[47]);
  FullAdder FA49 (Partial_Product[9][7],Partial_Product[10][6],Partial_Product[11][5],Sum[48],Carry_out[48]);
  FullAdder FA50 (Partial_Product[12][4],Partial_Product[13][3],Partial_Product[14][2],Sum[49],Carry_out[49]);
  HalfAdder HA51 (Partial_Product[15][1],Partial_Product[16][0],Sum[50],Carry_out[50]);
  FullAdder FA52 (Partial_Product[0][17],Partial_Product[1][16],Partial_Product[2][15],Sum[51],Carry_out[51]);
  FullAdder FA53 (Partial_Product[3][14],Partial_Product[4][13],Partial_Product[5][12],Sum[52],Carry_out[52]);
  FullAdder FA54 (Partial_Product[6][11],Partial_Product[7][10],Partial_Product[8][9],Sum[53],Carry_out[53]);
  FullAdder FA55 (Partial_Product[9][8],Partial_Product[10][7],Partial_Product[11][6],Sum[54],Carry_out[54]);
  FullAdder FA56 (Partial_Product[12][5],Partial_Product[13][4],Partial_Product[14][3],Sum[55],Carry_out[55]);
  FullAdder FA57 (Partial_Product[15][2],Partial_Product[16][1],Partial_Product[17][0],Sum[56],Carry_out[56]);
  FullAdder FA58 (Partial_Product[0][18],Partial_Product[1][17],Partial_Product[2][16],Sum[57],Carry_out[57]);
  FullAdder FA59 (Partial_Product[3][15],Partial_Product[4][14],Partial_Product[5][13],Sum[58],Carry_out[58]);
  FullAdder FA60 (Partial_Product[6][12],Partial_Product[7][11],Partial_Product[8][10],Sum[59],Carry_out[59]);
  FullAdder FA61 (Partial_Product[9][9],Partial_Product[10][8],Partial_Product[11][7],Sum[60],Carry_out[60]);
  FullAdder FA62 (Partial_Product[12][6],Partial_Product[13][5],Partial_Product[14][4],Sum[61],Carry_out[61]);
  FullAdder FA63 (Partial_Product[15][3],Partial_Product[16][2],Partial_Product[17][1],Sum[62],Carry_out[62]);
  FullAdder FA64 (Partial_Product[0][19],Partial_Product[1][18],Partial_Product[2][17],Sum[63],Carry_out[63]);
  FullAdder FA65 (Partial_Product[3][16],Partial_Product[4][15],Partial_Product[5][14],Sum[64],Carry_out[64]);
  FullAdder FA66 (Partial_Product[6][13],Partial_Product[7][12],Partial_Product[8][11],Sum[65],Carry_out[65]);
  FullAdder FA67 (Partial_Product[9][10],Partial_Product[10][9],Partial_Product[11][8],Sum[66],Carry_out[66]);
  FullAdder FA68 (Partial_Product[12][7],Partial_Product[13][6],Partial_Product[14][5],Sum[67],Carry_out[67]);
  FullAdder FA69 (Partial_Product[15][4],Partial_Product[16][3],Partial_Product[17][2],Sum[68],Carry_out[68]);
  HalfAdder HA70 (Partial_Product[18][1],Partial_Product[19][0],Sum[69],Carry_out[69]);
  FullAdder FA71 (Partial_Product[0][20],Partial_Product[1][19],Partial_Product[2][18],Sum[70],Carry_out[70]);
  FullAdder FA72 (Partial_Product[3][17],Partial_Product[4][16],Partial_Product[5][15],Sum[71],Carry_out[71]);
  FullAdder FA73 (Partial_Product[6][14],Partial_Product[7][13],Partial_Product[8][12],Sum[72],Carry_out[72]);
  FullAdder FA74 (Partial_Product[9][11],Partial_Product[10][10],Partial_Product[11][9],Sum[73],Carry_out[73]);
  FullAdder FA75 (Partial_Product[12][8],Partial_Product[13][7],Partial_Product[14][6],Sum[74],Carry_out[74]);
  FullAdder FA76 (Partial_Product[15][5],Partial_Product[16][4],Partial_Product[17][3],Sum[75],Carry_out[75]);
  FullAdder FA77 (Partial_Product[18][2],Partial_Product[19][1],Partial_Product[20][0],Sum[76],Carry_out[76]);
  FullAdder FA78 (Partial_Product[0][21],Partial_Product[1][20],Partial_Product[2][19],Sum[77],Carry_out[77]);
  FullAdder FA79 (Partial_Product[3][18],Partial_Product[4][17],Partial_Product[5][16],Sum[78],Carry_out[78]);
  FullAdder FA80 (Partial_Product[6][15],Partial_Product[7][14],Partial_Product[8][13],Sum[79],Carry_out[79]);
  FullAdder FA81 (Partial_Product[9][12],Partial_Product[10][11],Partial_Product[11][10],Sum[80],Carry_out[80]);
  FullAdder FA82 (Partial_Product[12][9],Partial_Product[13][8],Partial_Product[14][7],Sum[81],Carry_out[81]);
  FullAdder FA83 (Partial_Product[15][6],Partial_Product[16][5],Partial_Product[17][4],Sum[82],Carry_out[82]);
  FullAdder FA84 (Partial_Product[18][3],Partial_Product[19][2],Partial_Product[20][1],Sum[83],Carry_out[83]);
  FullAdder FA85 (Partial_Product[0][22],Partial_Product[1][21],Partial_Product[2][20],Sum[84],Carry_out[84]);
  FullAdder FA86 (Partial_Product[3][19],Partial_Product[4][18],Partial_Product[5][17],Sum[85],Carry_out[85]);
  FullAdder FA87 (Partial_Product[6][16],Partial_Product[7][15],Partial_Product[8][14],Sum[86],Carry_out[86]);
  FullAdder FA88 (Partial_Product[9][13],Partial_Product[10][12],Partial_Product[11][11],Sum[87],Carry_out[87]);
  FullAdder FA89 (Partial_Product[12][10],Partial_Product[13][9],Partial_Product[14][8],Sum[88],Carry_out[88]);
  FullAdder FA90 (Partial_Product[15][7],Partial_Product[16][6],Partial_Product[17][5],Sum[89],Carry_out[89]);
  FullAdder FA91 (Partial_Product[18][4],Partial_Product[19][3],Partial_Product[20][2],Sum[90],Carry_out[90]);
  HalfAdder HA92 (Partial_Product[21][1],Partial_Product[22][0],Sum[91],Carry_out[91]);
  FullAdder FA93 (Partial_Product[0][23],Partial_Product[1][22],Partial_Product[2][21],Sum[92],Carry_out[92]);
  FullAdder FA94 (Partial_Product[3][20],Partial_Product[4][19],Partial_Product[5][18],Sum[93],Carry_out[93]);
  FullAdder FA95 (Partial_Product[6][17],Partial_Product[7][16],Partial_Product[8][15],Sum[94],Carry_out[94]);
  FullAdder FA96 (Partial_Product[9][14],Partial_Product[10][13],Partial_Product[11][12],Sum[95],Carry_out[95]);
  FullAdder FA97 (Partial_Product[12][11],Partial_Product[13][10],Partial_Product[14][9],Sum[96],Carry_out[96]);
  FullAdder FA98 (Partial_Product[15][8],Partial_Product[16][7],Partial_Product[17][6],Sum[97],Carry_out[97]);
  FullAdder FA99 (Partial_Product[18][5],Partial_Product[19][4],Partial_Product[20][3],Sum[98],Carry_out[98]);
  FullAdder FA100 (Partial_Product[21][2],Partial_Product[22][1],Partial_Product[23][0],Sum[99],Carry_out[99]);
  FullAdder FA101 (Partial_Product[0][24],Partial_Product[1][23],Partial_Product[2][22],Sum[100],Carry_out[100]);
  FullAdder FA102 (Partial_Product[3][21],Partial_Product[4][20],Partial_Product[5][19],Sum[101],Carry_out[101]);
  FullAdder FA103 (Partial_Product[6][18],Partial_Product[7][17],Partial_Product[8][16],Sum[102],Carry_out[102]);
  FullAdder FA104 (Partial_Product[9][15],Partial_Product[10][14],Partial_Product[11][13],Sum[103],Carry_out[103]);
  FullAdder FA105 (Partial_Product[12][12],Partial_Product[13][11],Partial_Product[14][10],Sum[104],Carry_out[104]);
  FullAdder FA106 (Partial_Product[15][9],Partial_Product[16][8],Partial_Product[17][7],Sum[105],Carry_out[105]);
  FullAdder FA107 (Partial_Product[18][6],Partial_Product[19][5],Partial_Product[20][4],Sum[106],Carry_out[106]);
  FullAdder FA108 (Partial_Product[21][3],Partial_Product[22][2],Partial_Product[23][1],Sum[107],Carry_out[107]);
  FullAdder FA109 (Partial_Product[0][25],Partial_Product[1][24],Partial_Product[2][23],Sum[108],Carry_out[108]);
  FullAdder FA110 (Partial_Product[3][22],Partial_Product[4][21],Partial_Product[5][20],Sum[109],Carry_out[109]);
  FullAdder FA111 (Partial_Product[6][19],Partial_Product[7][18],Partial_Product[8][17],Sum[110],Carry_out[110]);
  FullAdder FA112 (Partial_Product[9][16],Partial_Product[10][15],Partial_Product[11][14],Sum[111],Carry_out[111]);
  FullAdder FA113 (Partial_Product[12][13],Partial_Product[13][12],Partial_Product[14][11],Sum[112],Carry_out[112]);
  FullAdder FA114 (Partial_Product[15][10],Partial_Product[16][9],Partial_Product[17][8],Sum[113],Carry_out[113]);
  FullAdder FA115 (Partial_Product[18][7],Partial_Product[19][6],Partial_Product[20][5],Sum[114],Carry_out[114]);
  FullAdder FA116 (Partial_Product[21][4],Partial_Product[22][3],Partial_Product[23][2],Sum[115],Carry_out[115]);
  HalfAdder HA117 (Partial_Product[24][1],Partial_Product[25][0],Sum[116],Carry_out[116]);
  FullAdder FA118 (Partial_Product[0][26],Partial_Product[1][25],Partial_Product[2][24],Sum[117],Carry_out[117]);
  FullAdder FA119 (Partial_Product[3][23],Partial_Product[4][22],Partial_Product[5][21],Sum[118],Carry_out[118]);
  FullAdder FA120 (Partial_Product[6][20],Partial_Product[7][19],Partial_Product[8][18],Sum[119],Carry_out[119]);
  FullAdder FA121 (Partial_Product[9][17],Partial_Product[10][16],Partial_Product[11][15],Sum[120],Carry_out[120]);
  FullAdder FA122 (Partial_Product[12][14],Partial_Product[13][13],Partial_Product[14][12],Sum[121],Carry_out[121]);
  FullAdder FA123 (Partial_Product[15][11],Partial_Product[16][10],Partial_Product[17][9],Sum[122],Carry_out[122]);
  FullAdder FA124 (Partial_Product[18][8],Partial_Product[19][7],Partial_Product[20][6],Sum[123],Carry_out[123]);
  FullAdder FA125 (Partial_Product[21][5],Partial_Product[22][4],Partial_Product[23][3],Sum[124],Carry_out[124]);
  FullAdder FA126 (Partial_Product[24][2],Partial_Product[25][1],Partial_Product[26][0],Sum[125],Carry_out[125]);
  FullAdder FA127 (Partial_Product[0][27],Partial_Product[1][26],Partial_Product[2][25],Sum[126],Carry_out[126]);
  FullAdder FA128 (Partial_Product[3][24],Partial_Product[4][23],Partial_Product[5][22],Sum[127],Carry_out[127]);
  FullAdder FA129 (Partial_Product[6][21],Partial_Product[7][20],Partial_Product[8][19],Sum[128],Carry_out[128]);
  FullAdder FA130 (Partial_Product[9][18],Partial_Product[10][17],Partial_Product[11][16],Sum[129],Carry_out[129]);
  FullAdder FA131 (Partial_Product[12][15],Partial_Product[13][14],Partial_Product[14][13],Sum[130],Carry_out[130]);
  FullAdder FA132 (Partial_Product[15][12],Partial_Product[16][11],Partial_Product[17][10],Sum[131],Carry_out[131]);
  FullAdder FA133 (Partial_Product[18][9],Partial_Product[19][8],Partial_Product[20][7],Sum[132],Carry_out[132]);
  FullAdder FA134 (Partial_Product[21][6],Partial_Product[22][5],Partial_Product[23][4],Sum[133],Carry_out[133]);
  FullAdder FA135 (Partial_Product[24][3],Partial_Product[25][2],Partial_Product[26][1],Sum[134],Carry_out[134]);
  FullAdder FA136 (Partial_Product[0][28],Partial_Product[1][27],Partial_Product[2][26],Sum[135],Carry_out[135]);
  FullAdder FA137 (Partial_Product[3][25],Partial_Product[4][24],Partial_Product[5][23],Sum[136],Carry_out[136]);
  FullAdder FA138 (Partial_Product[6][22],Partial_Product[7][21],Partial_Product[8][20],Sum[137],Carry_out[137]);
  FullAdder FA139 (Partial_Product[9][19],Partial_Product[10][18],Partial_Product[11][17],Sum[138],Carry_out[138]);
  FullAdder FA140 (Partial_Product[12][16],Partial_Product[13][15],Partial_Product[14][14],Sum[139],Carry_out[139]);
  FullAdder FA141 (Partial_Product[15][13],Partial_Product[16][12],Partial_Product[17][11],Sum[140],Carry_out[140]);
  FullAdder FA142 (Partial_Product[18][10],Partial_Product[19][9],Partial_Product[20][8],Sum[141],Carry_out[141]);
  FullAdder FA143 (Partial_Product[21][7],Partial_Product[22][6],Partial_Product[23][5],Sum[142],Carry_out[142]);
  FullAdder FA144 (Partial_Product[24][4],Partial_Product[25][3],Partial_Product[26][2],Sum[143],Carry_out[143]);
  HalfAdder HA145 (Partial_Product[27][1],Partial_Product[28][0],Sum[144],Carry_out[144]);
  FullAdder FA146 (Partial_Product[0][29],Partial_Product[1][28],Partial_Product[2][27],Sum[145],Carry_out[145]);
  FullAdder FA147 (Partial_Product[3][26],Partial_Product[4][25],Partial_Product[5][24],Sum[146],Carry_out[146]);
  FullAdder FA148 (Partial_Product[6][23],Partial_Product[7][22],Partial_Product[8][21],Sum[147],Carry_out[147]);
  FullAdder FA149 (Partial_Product[9][20],Partial_Product[10][19],Partial_Product[11][18],Sum[148],Carry_out[148]);
  FullAdder FA150 (Partial_Product[12][17],Partial_Product[13][16],Partial_Product[14][15],Sum[149],Carry_out[149]);
  FullAdder FA151 (Partial_Product[15][14],Partial_Product[16][13],Partial_Product[17][12],Sum[150],Carry_out[150]);
  FullAdder FA152 (Partial_Product[18][11],Partial_Product[19][10],Partial_Product[20][9],Sum[151],Carry_out[151]);
  FullAdder FA153 (Partial_Product[21][8],Partial_Product[22][7],Partial_Product[23][6],Sum[152],Carry_out[152]);
  FullAdder FA154 (Partial_Product[24][5],Partial_Product[25][4],Partial_Product[26][3],Sum[153],Carry_out[153]);
  FullAdder FA155 (Partial_Product[27][2],Partial_Product[28][1],Partial_Product[29][0],Sum[154],Carry_out[154]);
  FullAdder FA156 (Partial_Product[0][30],Partial_Product[1][29],Partial_Product[2][28],Sum[155],Carry_out[155]);
  FullAdder FA157 (Partial_Product[3][27],Partial_Product[4][26],Partial_Product[5][25],Sum[156],Carry_out[156]);
  FullAdder FA158 (Partial_Product[6][24],Partial_Product[7][23],Partial_Product[8][22],Sum[157],Carry_out[157]);
  FullAdder FA159 (Partial_Product[9][21],Partial_Product[10][20],Partial_Product[11][19],Sum[158],Carry_out[158]);
  FullAdder FA160 (Partial_Product[12][18],Partial_Product[13][17],Partial_Product[14][16],Sum[159],Carry_out[159]);
  FullAdder FA161 (Partial_Product[15][15],Partial_Product[16][14],Partial_Product[17][13],Sum[160],Carry_out[160]);
  FullAdder FA162 (Partial_Product[18][12],Partial_Product[19][11],Partial_Product[20][10],Sum[161],Carry_out[161]);
  FullAdder FA163 (Partial_Product[21][9],Partial_Product[22][8],Partial_Product[23][7],Sum[162],Carry_out[162]);
  FullAdder FA164 (Partial_Product[24][6],Partial_Product[25][5],Partial_Product[26][4],Sum[163],Carry_out[163]);
  FullAdder FA165 (Partial_Product[27][3],Partial_Product[28][2],Partial_Product[29][1],Sum[164],Carry_out[164]);
  FullAdder FA166 (Partial_Product[0][31],Partial_Product[1][30],Partial_Product[2][29],Sum[165],Carry_out[165]);
  FullAdder FA167 (Partial_Product[3][28],Partial_Product[4][27],Partial_Product[5][26],Sum[166],Carry_out[166]);
  FullAdder FA168 (Partial_Product[6][25],Partial_Product[7][24],Partial_Product[8][23],Sum[167],Carry_out[167]);
  FullAdder FA169 (Partial_Product[9][22],Partial_Product[10][21],Partial_Product[11][20],Sum[168],Carry_out[168]);
  FullAdder FA170 (Partial_Product[12][19],Partial_Product[13][18],Partial_Product[14][17],Sum[169],Carry_out[169]);
  FullAdder FA171 (Partial_Product[15][16],Partial_Product[16][15],Partial_Product[17][14],Sum[170],Carry_out[170]);
  FullAdder FA172 (Partial_Product[18][13],Partial_Product[19][12],Partial_Product[20][11],Sum[171],Carry_out[171]);
  FullAdder FA173 (Partial_Product[21][10],Partial_Product[22][9],Partial_Product[23][8],Sum[172],Carry_out[172]);
  FullAdder FA174 (Partial_Product[24][7],Partial_Product[25][6],Partial_Product[26][5],Sum[173],Carry_out[173]);
  FullAdder FA175 (Partial_Product[27][4],Partial_Product[28][3],Partial_Product[29][2],Sum[174],Carry_out[174]);
  FullAdder FA176 (Partial_Product[1][31],Partial_Product[2][30],Partial_Product[3][29],Sum[175],Carry_out[175]);
  FullAdder FA177 (Partial_Product[4][28],Partial_Product[5][27],Partial_Product[6][26],Sum[176],Carry_out[176]);
  FullAdder FA178 (Partial_Product[7][25],Partial_Product[8][24],Partial_Product[9][23],Sum[177],Carry_out[177]);
  FullAdder FA179 (Partial_Product[10][22],Partial_Product[11][21],Partial_Product[12][20],Sum[178],Carry_out[178]);
  FullAdder FA180 (Partial_Product[13][19],Partial_Product[14][18],Partial_Product[15][17],Sum[179],Carry_out[179]);
  FullAdder FA181 (Partial_Product[16][16],Partial_Product[17][15],Partial_Product[18][14],Sum[180],Carry_out[180]);
  FullAdder FA182 (Partial_Product[19][13],Partial_Product[20][12],Partial_Product[21][11],Sum[181],Carry_out[181]);
  FullAdder FA183 (Partial_Product[22][10],Partial_Product[23][9],Partial_Product[24][8],Sum[182],Carry_out[182]);
  FullAdder FA184 (Partial_Product[25][7],Partial_Product[26][6],Partial_Product[27][5],Sum[183],Carry_out[183]);
  HalfAdder HA185 (Partial_Product[28][4],Partial_Product[29][3],Sum[184],Carry_out[184]);
  FullAdder FA186 (Partial_Product[2][31],Partial_Product[3][30],Partial_Product[4][29],Sum[185],Carry_out[185]);
  FullAdder FA187 (Partial_Product[5][28],Partial_Product[6][27],Partial_Product[7][26],Sum[186],Carry_out[186]);
  FullAdder FA188 (Partial_Product[8][25],Partial_Product[9][24],Partial_Product[10][23],Sum[187],Carry_out[187]);
  FullAdder FA189 (Partial_Product[11][22],Partial_Product[12][21],Partial_Product[13][20],Sum[188],Carry_out[188]);
  FullAdder FA190 (Partial_Product[14][19],Partial_Product[15][18],Partial_Product[16][17],Sum[189],Carry_out[189]);
  FullAdder FA191 (Partial_Product[17][16],Partial_Product[18][15],Partial_Product[19][14],Sum[190],Carry_out[190]);
  FullAdder FA192 (Partial_Product[20][13],Partial_Product[21][12],Partial_Product[22][11],Sum[191],Carry_out[191]);
  FullAdder FA193 (Partial_Product[23][10],Partial_Product[24][9],Partial_Product[25][8],Sum[192],Carry_out[192]);
  FullAdder FA194 (Partial_Product[26][7],Partial_Product[27][6],Partial_Product[28][5],Sum[193],Carry_out[193]);
  FullAdder FA195 (Partial_Product[3][31],Partial_Product[4][30],Partial_Product[5][29],Sum[194],Carry_out[194]);
  FullAdder FA196 (Partial_Product[6][28],Partial_Product[7][27],Partial_Product[8][26],Sum[195],Carry_out[195]);
  FullAdder FA197 (Partial_Product[9][25],Partial_Product[10][24],Partial_Product[11][23],Sum[196],Carry_out[196]);
  FullAdder FA198 (Partial_Product[12][22],Partial_Product[13][21],Partial_Product[14][20],Sum[197],Carry_out[197]);
  FullAdder FA199 (Partial_Product[15][19],Partial_Product[16][18],Partial_Product[17][17],Sum[198],Carry_out[198]);
  FullAdder FA200 (Partial_Product[18][16],Partial_Product[19][15],Partial_Product[20][14],Sum[199],Carry_out[199]);
  FullAdder FA201 (Partial_Product[21][13],Partial_Product[22][12],Partial_Product[23][11],Sum[200],Carry_out[200]);
  FullAdder FA202 (Partial_Product[24][10],Partial_Product[25][9],Partial_Product[26][8],Sum[201],Carry_out[201]);
  FullAdder FA203 (Partial_Product[27][7],Partial_Product[28][6],Partial_Product[29][5],Sum[202],Carry_out[202]);
  FullAdder FA204 (Partial_Product[4][31],Partial_Product[5][30],Partial_Product[6][29],Sum[203],Carry_out[203]);
  FullAdder FA205 (Partial_Product[7][28],Partial_Product[8][27],Partial_Product[9][26],Sum[204],Carry_out[204]);
  FullAdder FA206 (Partial_Product[10][25],Partial_Product[11][24],Partial_Product[12][23],Sum[205],Carry_out[205]);
  FullAdder FA207 (Partial_Product[13][22],Partial_Product[14][21],Partial_Product[15][20],Sum[206],Carry_out[206]);
  FullAdder FA208 (Partial_Product[16][19],Partial_Product[17][18],Partial_Product[18][17],Sum[207],Carry_out[207]);
  FullAdder FA209 (Partial_Product[19][16],Partial_Product[20][15],Partial_Product[21][14],Sum[208],Carry_out[208]);
  FullAdder FA210 (Partial_Product[22][13],Partial_Product[23][12],Partial_Product[24][11],Sum[209],Carry_out[209]);
  FullAdder FA211 (Partial_Product[25][10],Partial_Product[26][9],Partial_Product[27][8],Sum[210],Carry_out[210]);
  HalfAdder HA212 (Partial_Product[28][7],Partial_Product[29][6],Sum[211],Carry_out[211]);
  FullAdder FA213 (Partial_Product[5][31],Partial_Product[6][30],Partial_Product[7][29],Sum[212],Carry_out[212]);
  FullAdder FA214 (Partial_Product[8][28],Partial_Product[9][27],Partial_Product[10][26],Sum[213],Carry_out[213]);
  FullAdder FA215 (Partial_Product[11][25],Partial_Product[12][24],Partial_Product[13][23],Sum[214],Carry_out[214]);
  FullAdder FA216 (Partial_Product[14][22],Partial_Product[15][21],Partial_Product[16][20],Sum[215],Carry_out[215]);
  FullAdder FA217 (Partial_Product[17][19],Partial_Product[18][18],Partial_Product[19][17],Sum[216],Carry_out[216]);
  FullAdder FA218 (Partial_Product[20][16],Partial_Product[21][15],Partial_Product[22][14],Sum[217],Carry_out[217]);
  FullAdder FA219 (Partial_Product[23][13],Partial_Product[24][12],Partial_Product[25][11],Sum[218],Carry_out[218]);
  FullAdder FA220 (Partial_Product[26][10],Partial_Product[27][9],Partial_Product[28][8],Sum[219],Carry_out[219]);
  FullAdder FA221 (Partial_Product[6][31],Partial_Product[7][30],Partial_Product[8][29],Sum[220],Carry_out[220]);
  FullAdder FA222 (Partial_Product[9][28],Partial_Product[10][27],Partial_Product[11][26],Sum[221],Carry_out[221]);
  FullAdder FA223 (Partial_Product[12][25],Partial_Product[13][24],Partial_Product[14][23],Sum[222],Carry_out[222]);
  FullAdder FA224 (Partial_Product[15][22],Partial_Product[16][21],Partial_Product[17][20],Sum[223],Carry_out[223]);
  FullAdder FA225 (Partial_Product[18][19],Partial_Product[19][18],Partial_Product[20][17],Sum[224],Carry_out[224]);
  FullAdder FA226 (Partial_Product[21][16],Partial_Product[22][15],Partial_Product[23][14],Sum[225],Carry_out[225]);
  FullAdder FA227 (Partial_Product[24][13],Partial_Product[25][12],Partial_Product[26][11],Sum[226],Carry_out[226]);
  FullAdder FA228 (Partial_Product[27][10],Partial_Product[28][9],Partial_Product[29][8],Sum[227],Carry_out[227]);
  FullAdder FA229 (Partial_Product[7][31],Partial_Product[8][30],Partial_Product[9][29],Sum[228],Carry_out[228]);
  FullAdder FA230 (Partial_Product[10][28],Partial_Product[11][27],Partial_Product[12][26],Sum[229],Carry_out[229]);
  FullAdder FA231 (Partial_Product[13][25],Partial_Product[14][24],Partial_Product[15][23],Sum[230],Carry_out[230]);
  FullAdder FA232 (Partial_Product[16][22],Partial_Product[17][21],Partial_Product[18][20],Sum[231],Carry_out[231]);
  FullAdder FA233 (Partial_Product[19][19],Partial_Product[20][18],Partial_Product[21][17],Sum[232],Carry_out[232]);
  FullAdder FA234 (Partial_Product[22][16],Partial_Product[23][15],Partial_Product[24][14],Sum[233],Carry_out[233]);
  FullAdder FA235 (Partial_Product[25][13],Partial_Product[26][12],Partial_Product[27][11],Sum[234],Carry_out[234]);
  HalfAdder HA236 (Partial_Product[28][10],Partial_Product[29][9],Sum[235],Carry_out[235]);
  FullAdder FA237 (Partial_Product[8][31],Partial_Product[9][30],Partial_Product[10][29],Sum[236],Carry_out[236]);
  FullAdder FA238 (Partial_Product[11][28],Partial_Product[12][27],Partial_Product[13][26],Sum[237],Carry_out[237]);
  FullAdder FA239 (Partial_Product[14][25],Partial_Product[15][24],Partial_Product[16][23],Sum[238],Carry_out[238]);
  FullAdder FA240 (Partial_Product[17][22],Partial_Product[18][21],Partial_Product[19][20],Sum[239],Carry_out[239]);
  FullAdder FA241 (Partial_Product[20][19],Partial_Product[21][18],Partial_Product[22][17],Sum[240],Carry_out[240]);
  FullAdder FA242 (Partial_Product[23][16],Partial_Product[24][15],Partial_Product[25][14],Sum[241],Carry_out[241]);
  FullAdder FA243 (Partial_Product[26][13],Partial_Product[27][12],Partial_Product[28][11],Sum[242],Carry_out[242]);
  FullAdder FA244 (Partial_Product[9][31],Partial_Product[10][30],Partial_Product[11][29],Sum[243],Carry_out[243]);
  FullAdder FA245 (Partial_Product[12][28],Partial_Product[13][27],Partial_Product[14][26],Sum[244],Carry_out[244]);
  FullAdder FA246 (Partial_Product[15][25],Partial_Product[16][24],Partial_Product[17][23],Sum[245],Carry_out[245]);
  FullAdder FA247 (Partial_Product[18][22],Partial_Product[19][21],Partial_Product[20][20],Sum[246],Carry_out[246]);
  FullAdder FA248 (Partial_Product[21][19],Partial_Product[22][18],Partial_Product[23][17],Sum[247],Carry_out[247]);
  FullAdder FA249 (Partial_Product[24][16],Partial_Product[25][15],Partial_Product[26][14],Sum[248],Carry_out[248]);
  FullAdder FA250 (Partial_Product[27][13],Partial_Product[28][12],Partial_Product[29][11],Sum[249],Carry_out[249]);
  FullAdder FA251 (Partial_Product[10][31],Partial_Product[11][30],Partial_Product[12][29],Sum[250],Carry_out[250]);
  FullAdder FA252 (Partial_Product[13][28],Partial_Product[14][27],Partial_Product[15][26],Sum[251],Carry_out[251]);
  FullAdder FA253 (Partial_Product[16][25],Partial_Product[17][24],Partial_Product[18][23],Sum[252],Carry_out[252]);
  FullAdder FA254 (Partial_Product[19][22],Partial_Product[20][21],Partial_Product[21][20],Sum[253],Carry_out[253]);
  FullAdder FA255 (Partial_Product[22][19],Partial_Product[23][18],Partial_Product[24][17],Sum[254],Carry_out[254]);
  FullAdder FA256 (Partial_Product[25][16],Partial_Product[26][15],Partial_Product[27][14],Sum[255],Carry_out[255]);
  HalfAdder HA257 (Partial_Product[28][13],Partial_Product[29][12],Sum[256],Carry_out[256]);
  FullAdder FA258 (Partial_Product[11][31],Partial_Product[12][30],Partial_Product[13][29],Sum[257],Carry_out[257]);
  FullAdder FA259 (Partial_Product[14][28],Partial_Product[15][27],Partial_Product[16][26],Sum[258],Carry_out[258]);
  FullAdder FA260 (Partial_Product[17][25],Partial_Product[18][24],Partial_Product[19][23],Sum[259],Carry_out[259]);
  FullAdder FA261 (Partial_Product[20][22],Partial_Product[21][21],Partial_Product[22][20],Sum[260],Carry_out[260]);
  FullAdder FA262 (Partial_Product[23][19],Partial_Product[24][18],Partial_Product[25][17],Sum[261],Carry_out[261]);
  FullAdder FA263 (Partial_Product[26][16],Partial_Product[27][15],Partial_Product[28][14],Sum[262],Carry_out[262]);
  FullAdder FA264 (Partial_Product[12][31],Partial_Product[13][30],Partial_Product[14][29],Sum[263],Carry_out[263]);
  FullAdder FA265 (Partial_Product[15][28],Partial_Product[16][27],Partial_Product[17][26],Sum[264],Carry_out[264]);
  FullAdder FA266 (Partial_Product[18][25],Partial_Product[19][24],Partial_Product[20][23],Sum[265],Carry_out[265]);
  FullAdder FA267 (Partial_Product[21][22],Partial_Product[22][21],Partial_Product[23][20],Sum[266],Carry_out[266]);
  FullAdder FA268 (Partial_Product[24][19],Partial_Product[25][18],Partial_Product[26][17],Sum[267],Carry_out[267]);
  FullAdder FA269 (Partial_Product[27][16],Partial_Product[28][15],Partial_Product[29][14],Sum[268],Carry_out[268]);
  FullAdder FA270 (Partial_Product[13][31],Partial_Product[14][30],Partial_Product[15][29],Sum[269],Carry_out[269]);
  FullAdder FA271 (Partial_Product[16][28],Partial_Product[17][27],Partial_Product[18][26],Sum[270],Carry_out[270]);
  FullAdder FA272 (Partial_Product[19][25],Partial_Product[20][24],Partial_Product[21][23],Sum[271],Carry_out[271]);
  FullAdder FA273 (Partial_Product[22][22],Partial_Product[23][21],Partial_Product[24][20],Sum[272],Carry_out[272]);
  FullAdder FA274 (Partial_Product[25][19],Partial_Product[26][18],Partial_Product[27][17],Sum[273],Carry_out[273]);
  HalfAdder HA275 (Partial_Product[28][16],Partial_Product[29][15],Sum[274],Carry_out[274]);
  FullAdder FA276 (Partial_Product[14][31],Partial_Product[15][30],Partial_Product[16][29],Sum[275],Carry_out[275]);
  FullAdder FA277 (Partial_Product[17][28],Partial_Product[18][27],Partial_Product[19][26],Sum[276],Carry_out[276]);
  FullAdder FA278 (Partial_Product[20][25],Partial_Product[21][24],Partial_Product[22][23],Sum[277],Carry_out[277]);
  FullAdder FA279 (Partial_Product[23][22],Partial_Product[24][21],Partial_Product[25][20],Sum[278],Carry_out[278]);
  FullAdder FA280 (Partial_Product[26][19],Partial_Product[27][18],Partial_Product[28][17],Sum[279],Carry_out[279]);
  FullAdder FA281 (Partial_Product[15][31],Partial_Product[16][30],Partial_Product[17][29],Sum[280],Carry_out[280]);
  FullAdder FA282 (Partial_Product[18][28],Partial_Product[19][27],Partial_Product[20][26],Sum[281],Carry_out[281]);
  FullAdder FA283 (Partial_Product[21][25],Partial_Product[22][24],Partial_Product[23][23],Sum[282],Carry_out[282]);
  FullAdder FA284 (Partial_Product[24][22],Partial_Product[25][21],Partial_Product[26][20],Sum[283],Carry_out[283]);
  FullAdder FA285 (Partial_Product[27][19],Partial_Product[28][18],Partial_Product[29][17],Sum[284],Carry_out[284]);
  FullAdder FA286 (Partial_Product[16][31],Partial_Product[17][30],Partial_Product[18][29],Sum[285],Carry_out[285]);
  FullAdder FA287 (Partial_Product[19][28],Partial_Product[20][27],Partial_Product[21][26],Sum[286],Carry_out[286]);
  FullAdder FA288 (Partial_Product[22][25],Partial_Product[23][24],Partial_Product[24][23],Sum[287],Carry_out[287]);
  FullAdder FA289 (Partial_Product[25][22],Partial_Product[26][21],Partial_Product[27][20],Sum[288],Carry_out[288]);
  HalfAdder HA290 (Partial_Product[28][19],Partial_Product[29][18],Sum[289],Carry_out[289]);
  FullAdder FA291 (Partial_Product[17][31],Partial_Product[18][30],Partial_Product[19][29],Sum[290],Carry_out[290]);
  FullAdder FA292 (Partial_Product[20][28],Partial_Product[21][27],Partial_Product[22][26],Sum[291],Carry_out[291]);
  FullAdder FA293 (Partial_Product[23][25],Partial_Product[24][24],Partial_Product[25][23],Sum[292],Carry_out[292]);
  FullAdder FA294 (Partial_Product[26][22],Partial_Product[27][21],Partial_Product[28][20],Sum[293],Carry_out[293]);
  FullAdder FA295 (Partial_Product[18][31],Partial_Product[19][30],Partial_Product[20][29],Sum[294],Carry_out[294]);
  FullAdder FA296 (Partial_Product[21][28],Partial_Product[22][27],Partial_Product[23][26],Sum[295],Carry_out[295]);
  FullAdder FA297 (Partial_Product[24][25],Partial_Product[25][24],Partial_Product[26][23],Sum[296],Carry_out[296]);
  FullAdder FA298 (Partial_Product[27][22],Partial_Product[28][21],Partial_Product[29][20],Sum[297],Carry_out[297]);
  FullAdder FA299 (Partial_Product[19][31],Partial_Product[20][30],Partial_Product[21][29],Sum[298],Carry_out[298]);
  FullAdder FA300 (Partial_Product[22][28],Partial_Product[23][27],Partial_Product[24][26],Sum[299],Carry_out[299]);
  FullAdder FA301 (Partial_Product[25][25],Partial_Product[26][24],Partial_Product[27][23],Sum[300],Carry_out[300]);
  HalfAdder HA302 (Partial_Product[28][22],Partial_Product[29][21],Sum[301],Carry_out[301]);
  FullAdder FA303 (Partial_Product[20][31],Partial_Product[21][30],Partial_Product[22][29],Sum[302],Carry_out[302]);
  FullAdder FA304 (Partial_Product[23][28],Partial_Product[24][27],Partial_Product[25][26],Sum[303],Carry_out[303]);
  FullAdder FA305 (Partial_Product[26][25],Partial_Product[27][24],Partial_Product[28][23],Sum[304],Carry_out[304]);
  FullAdder FA306 (Partial_Product[21][31],Partial_Product[22][30],Partial_Product[23][29],Sum[305],Carry_out[305]);
  FullAdder FA307 (Partial_Product[24][28],Partial_Product[25][27],Partial_Product[26][26],Sum[306],Carry_out[306]);
  FullAdder FA308 (Partial_Product[27][25],Partial_Product[28][24],Partial_Product[29][23],Sum[307],Carry_out[307]);
  FullAdder FA309 (Partial_Product[22][31],Partial_Product[23][30],Partial_Product[24][29],Sum[308],Carry_out[308]);
  FullAdder FA310 (Partial_Product[25][28],Partial_Product[26][27],Partial_Product[27][26],Sum[309],Carry_out[309]);
  HalfAdder HA311 (Partial_Product[28][25],Partial_Product[29][24],Sum[310],Carry_out[310]);
  FullAdder FA312 (Partial_Product[23][31],Partial_Product[24][30],Partial_Product[25][29],Sum[311],Carry_out[311]);
  FullAdder FA313 (Partial_Product[26][28],Partial_Product[27][27],Partial_Product[28][26],Sum[312],Carry_out[312]);
  FullAdder FA314 (Partial_Product[24][31],Partial_Product[25][30],Partial_Product[26][29],Sum[313],Carry_out[313]);
  FullAdder FA315 (Partial_Product[27][28],Partial_Product[28][27],Partial_Product[29][26],Sum[314],Carry_out[314]);
  FullAdder FA316 (Partial_Product[25][31],Partial_Product[26][30],Partial_Product[27][29],Sum[315],Carry_out[315]);
  HalfAdder HA317 (Partial_Product[28][28],Partial_Product[29][27],Sum[316],Carry_out[316]);
  FullAdder FA318 (Partial_Product[26][31],Partial_Product[27][30],Partial_Product[28][29],Sum[317],Carry_out[317]);
  FullAdder FA319 (Partial_Product[27][31],Partial_Product[28][30],Partial_Product[29][29],Sum[318],Carry_out[318]);
  HalfAdder HA320 (Partial_Product[28][31],Partial_Product[29][30],Sum[319],Carry_out[319]);
  HalfAdder HA321 (Carry_out[0],Sum[1],Sum[320],Carry_out[320]);
  FullAdder FA322 (Partial_Product[3][0],Carry_out[1],Sum[2],Sum[321],Carry_out[321]);
  FullAdder FA323 (Carry_out[2],Sum[3],Sum[4],Sum[322],Carry_out[322]);
  FullAdder FA324 (Carry_out[3],Carry_out[4],Sum[5],Sum[323],Carry_out[323]);
  FullAdder FA325 (Partial_Product[6][0],Carry_out[5],Carry_out[6],Sum[324],Carry_out[324]);
  HalfAdder HA326 (Sum[7],Sum[8],Sum[325],Carry_out[325]);
  FullAdder FA327 (Carry_out[7],Carry_out[8],Sum[9],Sum[326],Carry_out[326]);
  HalfAdder HA328 (Sum[10],Sum[11],Sum[327],Carry_out[327]);
  FullAdder FA329 (Carry_out[9],Carry_out[10],Carry_out[11],Sum[328],Carry_out[328]);
  FullAdder FA330 (Sum[12],Sum[13],Sum[14],Sum[329],Carry_out[329]);
  FullAdder FA331 (Partial_Product[9][0],Carry_out[12],Carry_out[13],Sum[330],Carry_out[330]);
  FullAdder FA332 (Carry_out[14],Sum[15],Sum[16],Sum[331],Carry_out[331]);
  FullAdder FA333 (Carry_out[15],Carry_out[16],Carry_out[17],Sum[332],Carry_out[332]);
  FullAdder FA334 (Sum[18],Sum[19],Sum[20],Sum[333],Carry_out[333]);
  FullAdder FA335 (Carry_out[18],Carry_out[19],Carry_out[20],Sum[334],Carry_out[334]);
  FullAdder FA336 (Carry_out[21],Sum[22],Sum[23],Sum[335],Carry_out[335]);
  HalfAdder HA337 (Sum[24],Sum[25],Sum[336],Carry_out[336]);
  FullAdder FA338 (Partial_Product[12][0],Carry_out[22],Carry_out[23],Sum[337],Carry_out[337]);
  FullAdder FA339 (Carry_out[24],Carry_out[25],Sum[26],Sum[338],Carry_out[338]);
  FullAdder FA340 (Sum[27],Sum[28],Sum[29],Sum[339],Carry_out[339]);
  FullAdder FA341 (Carry_out[26],Carry_out[27],Carry_out[28],Sum[340],Carry_out[340]);
  FullAdder FA342 (Carry_out[29],Sum[30],Sum[31],Sum[341],Carry_out[341]);
  FullAdder FA343 (Sum[32],Sum[33],Sum[34],Sum[342],Carry_out[342]);
  FullAdder FA344 (Carry_out[30],Carry_out[31],Carry_out[32],Sum[343],Carry_out[343]);
  FullAdder FA345 (Carry_out[33],Carry_out[34],Sum[35],Sum[344],Carry_out[344]);
  FullAdder FA346 (Sum[36],Sum[37],Sum[38],Sum[345],Carry_out[345]);
  FullAdder FA347 (Partial_Product[15][0],Carry_out[35],Carry_out[36],Sum[346],Carry_out[346]);
  FullAdder FA348 (Carry_out[37],Carry_out[38],Carry_out[39],Sum[347],Carry_out[347]);
  FullAdder FA349 (Sum[40],Sum[41],Sum[42],Sum[348],Carry_out[348]);
  HalfAdder HA350 (Sum[43],Sum[44],Sum[349],Carry_out[349]);
  FullAdder FA351 (Carry_out[40],Carry_out[41],Carry_out[42],Sum[350],Carry_out[350]);
  FullAdder FA352 (Carry_out[43],Carry_out[44],Sum[45],Sum[351],Carry_out[351]);
  FullAdder FA353 (Sum[46],Sum[47],Sum[48],Sum[352],Carry_out[352]);
  HalfAdder HA354 (Sum[49],Sum[50],Sum[353],Carry_out[353]);
  FullAdder FA355 (Carry_out[45],Carry_out[46],Carry_out[47],Sum[354],Carry_out[354]);
  FullAdder FA356 (Carry_out[48],Carry_out[49],Carry_out[50],Sum[355],Carry_out[355]);
  FullAdder FA357 (Sum[51],Sum[52],Sum[53],Sum[356],Carry_out[356]);
  FullAdder FA358 (Sum[54],Sum[55],Sum[56],Sum[357],Carry_out[357]);
  FullAdder FA359 (Partial_Product[18][0],Carry_out[51],Carry_out[52],Sum[358],Carry_out[358]);
  FullAdder FA360 (Carry_out[53],Carry_out[54],Carry_out[55],Sum[359],Carry_out[359]);
  FullAdder FA361 (Carry_out[56],Sum[57],Sum[58],Sum[360],Carry_out[360]);
  FullAdder FA362 (Sum[59],Sum[60],Sum[61],Sum[361],Carry_out[361]);
  FullAdder FA363 (Carry_out[57],Carry_out[58],Carry_out[59],Sum[362],Carry_out[362]);
  FullAdder FA364 (Carry_out[60],Carry_out[61],Carry_out[62],Sum[363],Carry_out[363]);
  FullAdder FA365 (Sum[63],Sum[64],Sum[65],Sum[364],Carry_out[364]);
  FullAdder FA366 (Sum[66],Sum[67],Sum[68],Sum[365],Carry_out[365]);
  FullAdder FA367 (Carry_out[63],Carry_out[64],Carry_out[65],Sum[366],Carry_out[366]);
  FullAdder FA368 (Carry_out[66],Carry_out[67],Carry_out[68],Sum[367],Carry_out[367]);
  FullAdder FA369 (Carry_out[69],Sum[70],Sum[71],Sum[368],Carry_out[368]);
  FullAdder FA370 (Sum[72],Sum[73],Sum[74],Sum[369],Carry_out[369]);
  HalfAdder HA371 (Sum[75],Sum[76],Sum[370],Carry_out[370]);
  FullAdder FA372 (Partial_Product[21][0],Carry_out[70],Carry_out[71],Sum[371],Carry_out[371]);
  FullAdder FA373 (Carry_out[72],Carry_out[73],Carry_out[74],Sum[372],Carry_out[372]);
  FullAdder FA374 (Carry_out[75],Carry_out[76],Sum[77],Sum[373],Carry_out[373]);
  FullAdder FA375 (Sum[78],Sum[79],Sum[80],Sum[374],Carry_out[374]);
  FullAdder FA376 (Sum[81],Sum[82],Sum[83],Sum[375],Carry_out[375]);
  FullAdder FA377 (Carry_out[77],Carry_out[78],Carry_out[79],Sum[376],Carry_out[376]);
  FullAdder FA378 (Carry_out[80],Carry_out[81],Carry_out[82],Sum[377],Carry_out[377]);
  FullAdder FA379 (Carry_out[83],Sum[84],Sum[85],Sum[378],Carry_out[378]);
  FullAdder FA380 (Sum[86],Sum[87],Sum[88],Sum[379],Carry_out[379]);
  FullAdder FA381 (Sum[89],Sum[90],Sum[91],Sum[380],Carry_out[380]);
  FullAdder FA382 (Carry_out[84],Carry_out[85],Carry_out[86],Sum[381],Carry_out[381]);
  FullAdder FA383 (Carry_out[87],Carry_out[88],Carry_out[89],Sum[382],Carry_out[382]);
  FullAdder FA384 (Carry_out[90],Carry_out[91],Sum[92],Sum[383],Carry_out[383]);
  FullAdder FA385 (Sum[93],Sum[94],Sum[95],Sum[384],Carry_out[384]);
  FullAdder FA386 (Sum[96],Sum[97],Sum[98],Sum[385],Carry_out[385]);
  FullAdder FA387 (Partial_Product[24][0],Carry_out[92],Carry_out[93],Sum[386],Carry_out[386]);
  FullAdder FA388 (Carry_out[94],Carry_out[95],Carry_out[96],Sum[387],Carry_out[387]);
  FullAdder FA389 (Carry_out[97],Carry_out[98],Carry_out[99],Sum[388],Carry_out[388]);
  FullAdder FA390 (Sum[100],Sum[101],Sum[102],Sum[389],Carry_out[389]);
  FullAdder FA391 (Sum[103],Sum[104],Sum[105],Sum[390],Carry_out[390]);
  HalfAdder HA392 (Sum[106],Sum[107],Sum[391],Carry_out[391]);
  FullAdder FA393 (Carry_out[100],Carry_out[101],Carry_out[102],Sum[392],Carry_out[392]);
  FullAdder FA394 (Carry_out[103],Carry_out[104],Carry_out[105],Sum[393],Carry_out[393]);
  FullAdder FA395 (Carry_out[106],Carry_out[107],Sum[108],Sum[394],Carry_out[394]);
  FullAdder FA396 (Sum[109],Sum[110],Sum[111],Sum[395],Carry_out[395]);
  FullAdder FA397 (Sum[112],Sum[113],Sum[114],Sum[396],Carry_out[396]);
  HalfAdder HA398 (Sum[115],Sum[116],Sum[397],Carry_out[397]);
  FullAdder FA399 (Carry_out[108],Carry_out[109],Carry_out[110],Sum[398],Carry_out[398]);
  FullAdder FA400 (Carry_out[111],Carry_out[112],Carry_out[113],Sum[399],Carry_out[399]);
  FullAdder FA401 (Carry_out[114],Carry_out[115],Carry_out[116],Sum[400],Carry_out[400]);
  FullAdder FA402 (Sum[117],Sum[118],Sum[119],Sum[401],Carry_out[401]);
  FullAdder FA403 (Sum[120],Sum[121],Sum[122],Sum[402],Carry_out[402]);
  FullAdder FA404 (Sum[123],Sum[124],Sum[125],Sum[403],Carry_out[403]);
  FullAdder FA405 (Partial_Product[27][0],Carry_out[117],Carry_out[118],Sum[404],Carry_out[404]);
  FullAdder FA406 (Carry_out[119],Carry_out[120],Carry_out[121],Sum[405],Carry_out[405]);
  FullAdder FA407 (Carry_out[122],Carry_out[123],Carry_out[124],Sum[406],Carry_out[406]);
  FullAdder FA408 (Carry_out[125],Sum[126],Sum[127],Sum[407],Carry_out[407]);
  FullAdder FA409 (Sum[128],Sum[129],Sum[130],Sum[408],Carry_out[408]);
  FullAdder FA410 (Sum[131],Sum[132],Sum[133],Sum[409],Carry_out[409]);
  FullAdder FA411 (Carry_out[126],Carry_out[127],Carry_out[128],Sum[410],Carry_out[410]);
  FullAdder FA412 (Carry_out[129],Carry_out[130],Carry_out[131],Sum[411],Carry_out[411]);
  FullAdder FA413 (Carry_out[132],Carry_out[133],Carry_out[134],Sum[412],Carry_out[412]);
  FullAdder FA414 (Sum[135],Sum[136],Sum[137],Sum[413],Carry_out[413]);
  FullAdder FA415 (Sum[138],Sum[139],Sum[140],Sum[414],Carry_out[414]);
  FullAdder FA416 (Sum[141],Sum[142],Sum[143],Sum[415],Carry_out[415]);
  FullAdder FA417 (Carry_out[135],Carry_out[136],Carry_out[137],Sum[416],Carry_out[416]);
  FullAdder FA418 (Carry_out[138],Carry_out[139],Carry_out[140],Sum[417],Carry_out[417]);
  FullAdder FA419 (Carry_out[141],Carry_out[142],Carry_out[143],Sum[418],Carry_out[418]);
  FullAdder FA420 (Carry_out[144],Sum[145],Sum[146],Sum[419],Carry_out[419]);
  FullAdder FA421 (Sum[147],Sum[148],Sum[149],Sum[420],Carry_out[420]);
  FullAdder FA422 (Sum[150],Sum[151],Sum[152],Sum[421],Carry_out[421]);
  HalfAdder HA423 (Sum[153],Sum[154],Sum[422],Carry_out[422]);
  FullAdder FA424 (Partial_Product[30][0],Carry_out[145],Carry_out[146],Sum[423],Carry_out[423]);
  FullAdder FA425 (Carry_out[147],Carry_out[148],Carry_out[149],Sum[424],Carry_out[424]);
  FullAdder FA426 (Carry_out[150],Carry_out[151],Carry_out[152],Sum[425],Carry_out[425]);
  FullAdder FA427 (Carry_out[153],Carry_out[154],Sum[155],Sum[426],Carry_out[426]);
  FullAdder FA428 (Sum[156],Sum[157],Sum[158],Sum[427],Carry_out[427]);
  FullAdder FA429 (Sum[159],Sum[160],Sum[161],Sum[428],Carry_out[428]);
  FullAdder FA430 (Sum[162],Sum[163],Sum[164],Sum[429],Carry_out[429]);
  FullAdder FA431 (Partial_Product[30][1],Partial_Product[31][0],Carry_out[155],Sum[430],Carry_out[430]);
  FullAdder FA432 (Carry_out[156],Carry_out[157],Carry_out[158],Sum[431],Carry_out[431]);
  FullAdder FA433 (Carry_out[159],Carry_out[160],Carry_out[161],Sum[432],Carry_out[432]);
  FullAdder FA434 (Carry_out[162],Carry_out[163],Carry_out[164],Sum[433],Carry_out[433]);
  FullAdder FA435 (Sum[165],Sum[166],Sum[167],Sum[434],Carry_out[434]);
  FullAdder FA436 (Sum[168],Sum[169],Sum[170],Sum[435],Carry_out[435]);
  FullAdder FA437 (Sum[171],Sum[172],Sum[173],Sum[436],Carry_out[436]);
  FullAdder FA438 (Partial_Product[30][2],Partial_Product[31][1],Carry_out[165],Sum[437],Carry_out[437]);
  FullAdder FA439 (Carry_out[166],Carry_out[167],Carry_out[168],Sum[438],Carry_out[438]);
  FullAdder FA440 (Carry_out[169],Carry_out[170],Carry_out[171],Sum[439],Carry_out[439]);
  FullAdder FA441 (Carry_out[172],Carry_out[173],Carry_out[174],Sum[440],Carry_out[440]);
  FullAdder FA442 (Sum[175],Sum[176],Sum[177],Sum[441],Carry_out[441]);
  FullAdder FA443 (Sum[178],Sum[179],Sum[180],Sum[442],Carry_out[442]);
  FullAdder FA444 (Sum[181],Sum[182],Sum[183],Sum[443],Carry_out[443]);
  FullAdder FA445 (Partial_Product[29][4],Partial_Product[30][3],Partial_Product[31][2],Sum[444],Carry_out[444]);
  FullAdder FA446 (Carry_out[175],Carry_out[176],Carry_out[177],Sum[445],Carry_out[445]);
  FullAdder FA447 (Carry_out[178],Carry_out[179],Carry_out[180],Sum[446],Carry_out[446]);
  FullAdder FA448 (Carry_out[181],Carry_out[182],Carry_out[183],Sum[447],Carry_out[447]);
  FullAdder FA449 (Carry_out[184],Sum[185],Sum[186],Sum[448],Carry_out[448]);
  FullAdder FA450 (Sum[187],Sum[188],Sum[189],Sum[449],Carry_out[449]);
  FullAdder FA451 (Sum[190],Sum[191],Sum[192],Sum[450],Carry_out[450]);
  FullAdder FA452 (Partial_Product[30][4],Partial_Product[31][3],Carry_out[185],Sum[451],Carry_out[451]);
  FullAdder FA453 (Carry_out[186],Carry_out[187],Carry_out[188],Sum[452],Carry_out[452]);
  FullAdder FA454 (Carry_out[189],Carry_out[190],Carry_out[191],Sum[453],Carry_out[453]);
  FullAdder FA455 (Carry_out[192],Carry_out[193],Sum[194],Sum[454],Carry_out[454]);
  FullAdder FA456 (Sum[195],Sum[196],Sum[197],Sum[455],Carry_out[455]);
  FullAdder FA457 (Sum[198],Sum[199],Sum[200],Sum[456],Carry_out[456]);
  FullAdder FA458 (Partial_Product[30][5],Partial_Product[31][4],Carry_out[194],Sum[457],Carry_out[457]);
  FullAdder FA459 (Carry_out[195],Carry_out[196],Carry_out[197],Sum[458],Carry_out[458]);
  FullAdder FA460 (Carry_out[198],Carry_out[199],Carry_out[200],Sum[459],Carry_out[459]);
  FullAdder FA461 (Carry_out[201],Carry_out[202],Sum[203],Sum[460],Carry_out[460]);
  FullAdder FA462 (Sum[204],Sum[205],Sum[206],Sum[461],Carry_out[461]);
  FullAdder FA463 (Sum[207],Sum[208],Sum[209],Sum[462],Carry_out[462]);
  FullAdder FA464 (Partial_Product[29][7],Partial_Product[30][6],Partial_Product[31][5],Sum[463],Carry_out[463]);
  FullAdder FA465 (Carry_out[203],Carry_out[204],Carry_out[205],Sum[464],Carry_out[464]);
  FullAdder FA466 (Carry_out[206],Carry_out[207],Carry_out[208],Sum[465],Carry_out[465]);
  FullAdder FA467 (Carry_out[209],Carry_out[210],Carry_out[211],Sum[466],Carry_out[466]);
  FullAdder FA468 (Sum[212],Sum[213],Sum[214],Sum[467],Carry_out[467]);
  FullAdder FA469 (Sum[215],Sum[216],Sum[217],Sum[468],Carry_out[468]);
  FullAdder FA470 (Partial_Product[30][7],Partial_Product[31][6],Carry_out[212],Sum[469],Carry_out[469]);
  FullAdder FA471 (Carry_out[213],Carry_out[214],Carry_out[215],Sum[470],Carry_out[470]);
  FullAdder FA472 (Carry_out[216],Carry_out[217],Carry_out[218],Sum[471],Carry_out[471]);
  FullAdder FA473 (Carry_out[219],Sum[220],Sum[221],Sum[472],Carry_out[472]);
  FullAdder FA474 (Sum[222],Sum[223],Sum[224],Sum[473],Carry_out[473]);
  HalfAdder HA475 (Sum[225],Sum[226],Sum[474],Carry_out[474]);
  FullAdder FA476 (Partial_Product[30][8],Partial_Product[31][7],Carry_out[220],Sum[475],Carry_out[475]);
  FullAdder FA477 (Carry_out[221],Carry_out[222],Carry_out[223],Sum[476],Carry_out[476]);
  FullAdder FA478 (Carry_out[224],Carry_out[225],Carry_out[226],Sum[477],Carry_out[477]);
  FullAdder FA479 (Carry_out[227],Sum[228],Sum[229],Sum[478],Carry_out[478]);
  FullAdder FA480 (Sum[230],Sum[231],Sum[232],Sum[479],Carry_out[479]);
  HalfAdder HA481 (Sum[233],Sum[234],Sum[480],Carry_out[480]);
  FullAdder FA482 (Partial_Product[29][10],Partial_Product[30][9],Partial_Product[31][8],Sum[481],Carry_out[481]);
  FullAdder FA483 (Carry_out[228],Carry_out[229],Carry_out[230],Sum[482],Carry_out[482]);
  FullAdder FA484 (Carry_out[231],Carry_out[232],Carry_out[233],Sum[483],Carry_out[483]);
  FullAdder FA485 (Carry_out[234],Carry_out[235],Sum[236],Sum[484],Carry_out[484]);
  FullAdder FA486 (Sum[237],Sum[238],Sum[239],Sum[485],Carry_out[485]);
  HalfAdder HA487 (Sum[240],Sum[241],Sum[486],Carry_out[486]);
  FullAdder FA488 (Partial_Product[30][10],Partial_Product[31][9],Carry_out[236],Sum[487],Carry_out[487]);
  FullAdder FA489 (Carry_out[237],Carry_out[238],Carry_out[239],Sum[488],Carry_out[488]);
  FullAdder FA490 (Carry_out[240],Carry_out[241],Carry_out[242],Sum[489],Carry_out[489]);
  FullAdder FA491 (Sum[243],Sum[244],Sum[245],Sum[490],Carry_out[490]);
  FullAdder FA492 (Sum[246],Sum[247],Sum[248],Sum[491],Carry_out[491]);
  FullAdder FA493 (Partial_Product[30][11],Partial_Product[31][10],Carry_out[243],Sum[492],Carry_out[492]);
  FullAdder FA494 (Carry_out[244],Carry_out[245],Carry_out[246],Sum[493],Carry_out[493]);
  FullAdder FA495 (Carry_out[247],Carry_out[248],Carry_out[249],Sum[494],Carry_out[494]);
  FullAdder FA496 (Sum[250],Sum[251],Sum[252],Sum[495],Carry_out[495]);
  FullAdder FA497 (Sum[253],Sum[254],Sum[255],Sum[496],Carry_out[496]);
  FullAdder FA498 (Partial_Product[29][13],Partial_Product[30][12],Partial_Product[31][11],Sum[497],Carry_out[497]);
  FullAdder FA499 (Carry_out[250],Carry_out[251],Carry_out[252],Sum[498],Carry_out[498]);
  FullAdder FA500 (Carry_out[253],Carry_out[254],Carry_out[255],Sum[499],Carry_out[499]);
  FullAdder FA501 (Carry_out[256],Sum[257],Sum[258],Sum[500],Carry_out[500]);
  FullAdder FA502 (Sum[259],Sum[260],Sum[261],Sum[501],Carry_out[501]);
  FullAdder FA503 (Partial_Product[30][13],Partial_Product[31][12],Carry_out[257],Sum[502],Carry_out[502]);
  FullAdder FA504 (Carry_out[258],Carry_out[259],Carry_out[260],Sum[503],Carry_out[503]);
  FullAdder FA505 (Carry_out[261],Carry_out[262],Sum[263],Sum[504],Carry_out[504]);
  FullAdder FA506 (Sum[264],Sum[265],Sum[266],Sum[505],Carry_out[505]);
  FullAdder FA507 (Partial_Product[30][14],Partial_Product[31][13],Carry_out[263],Sum[506],Carry_out[506]);
  FullAdder FA508 (Carry_out[264],Carry_out[265],Carry_out[266],Sum[507],Carry_out[507]);
  FullAdder FA509 (Carry_out[267],Carry_out[268],Sum[269],Sum[508],Carry_out[508]);
  FullAdder FA510 (Sum[270],Sum[271],Sum[272],Sum[509],Carry_out[509]);
  FullAdder FA511 (Partial_Product[29][16],Partial_Product[30][15],Partial_Product[31][14],Sum[510],Carry_out[510]);
  FullAdder FA512 (Carry_out[269],Carry_out[270],Carry_out[271],Sum[511],Carry_out[511]);
  FullAdder FA513 (Carry_out[272],Carry_out[273],Carry_out[274],Sum[512],Carry_out[512]);
  FullAdder FA514 (Sum[275],Sum[276],Sum[277],Sum[513],Carry_out[513]);
  FullAdder FA515 (Partial_Product[30][16],Partial_Product[31][15],Carry_out[275],Sum[514],Carry_out[514]);
  FullAdder FA516 (Carry_out[276],Carry_out[277],Carry_out[278],Sum[515],Carry_out[515]);
  FullAdder FA517 (Carry_out[279],Sum[280],Sum[281],Sum[516],Carry_out[516]);
  HalfAdder HA518 (Sum[282],Sum[283],Sum[517],Carry_out[517]);
  FullAdder FA519 (Partial_Product[30][17],Partial_Product[31][16],Carry_out[280],Sum[518],Carry_out[518]);
  FullAdder FA520 (Carry_out[281],Carry_out[282],Carry_out[283],Sum[519],Carry_out[519]);
  FullAdder FA521 (Carry_out[284],Sum[285],Sum[286],Sum[520],Carry_out[520]);
  HalfAdder HA522 (Sum[287],Sum[288],Sum[521],Carry_out[521]);
  FullAdder FA523 (Partial_Product[29][19],Partial_Product[30][18],Partial_Product[31][17],Sum[522],Carry_out[522]);
  FullAdder FA524 (Carry_out[285],Carry_out[286],Carry_out[287],Sum[523],Carry_out[523]);
  FullAdder FA525 (Carry_out[288],Carry_out[289],Sum[290],Sum[524],Carry_out[524]);
  HalfAdder HA526 (Sum[291],Sum[292],Sum[525],Carry_out[525]);
  FullAdder FA527 (Partial_Product[30][19],Partial_Product[31][18],Carry_out[290],Sum[526],Carry_out[526]);
  FullAdder FA528 (Carry_out[291],Carry_out[292],Carry_out[293],Sum[527],Carry_out[527]);
  FullAdder FA529 (Sum[294],Sum[295],Sum[296],Sum[528],Carry_out[528]);
  FullAdder FA530 (Partial_Product[30][20],Partial_Product[31][19],Carry_out[294],Sum[529],Carry_out[529]);
  FullAdder FA531 (Carry_out[295],Carry_out[296],Carry_out[297],Sum[530],Carry_out[530]);
  FullAdder FA532 (Sum[298],Sum[299],Sum[300],Sum[531],Carry_out[531]);
  FullAdder FA533 (Partial_Product[29][22],Partial_Product[30][21],Partial_Product[31][20],Sum[532],Carry_out[532]);
  FullAdder FA534 (Carry_out[298],Carry_out[299],Carry_out[300],Sum[533],Carry_out[533]);
  FullAdder FA535 (Carry_out[301],Sum[302],Sum[303],Sum[534],Carry_out[534]);
  FullAdder FA536 (Partial_Product[30][22],Partial_Product[31][21],Carry_out[302],Sum[535],Carry_out[535]);
  FullAdder FA537 (Carry_out[303],Carry_out[304],Sum[305],Sum[536],Carry_out[536]);
  FullAdder FA538 (Partial_Product[30][23],Partial_Product[31][22],Carry_out[305],Sum[537],Carry_out[537]);
  FullAdder FA539 (Carry_out[306],Carry_out[307],Sum[308],Sum[538],Carry_out[538]);
  FullAdder FA540 (Partial_Product[29][25],Partial_Product[30][24],Partial_Product[31][23],Sum[539],Carry_out[539]);
  FullAdder FA541 (Carry_out[308],Carry_out[309],Carry_out[310],Sum[540],Carry_out[540]);
  FullAdder FA542 (Partial_Product[30][25],Partial_Product[31][24],Carry_out[311],Sum[541],Carry_out[541]);
  HalfAdder HA543 (Carry_out[312],Sum[313],Sum[542],Carry_out[542]);
  FullAdder FA544 (Partial_Product[30][26],Partial_Product[31][25],Carry_out[313],Sum[543],Carry_out[543]);
  HalfAdder HA545 (Carry_out[314],Sum[315],Sum[544],Carry_out[544]);
  FullAdder FA546 (Partial_Product[29][28],Partial_Product[30][27],Partial_Product[31][26],Sum[545],Carry_out[545]);
  HalfAdder HA547 (Carry_out[315],Carry_out[316],Sum[546],Carry_out[546]);
  FullAdder FA548 (Partial_Product[30][28],Partial_Product[31][27],Carry_out[317],Sum[547],Carry_out[547]);
  FullAdder FA549 (Partial_Product[30][29],Partial_Product[31][28],Carry_out[318],Sum[548],Carry_out[548]);
  FullAdder FA550 (Partial_Product[29][31],Partial_Product[30][30],Partial_Product[31][29],Sum[549],Carry_out[549]);
  HalfAdder HA551 (Carry_out[320],Sum[321],Sum[550],Carry_out[550]);
  HalfAdder HA552 (Carry_out[321],Sum[322],Sum[551],Carry_out[551]);
  FullAdder FA553 (Sum[6],Carry_out[322],Sum[323],Sum[552],Carry_out[552]);
  FullAdder FA554 (Carry_out[323],Sum[324],Sum[325],Sum[553],Carry_out[553]);
  FullAdder FA555 (Carry_out[324],Carry_out[325],Sum[326],Sum[554],Carry_out[554]);
  FullAdder FA556 (Carry_out[326],Carry_out[327],Sum[328],Sum[555],Carry_out[555]);
  FullAdder FA557 (Sum[17],Carry_out[328],Carry_out[329],Sum[556],Carry_out[556]);
  HalfAdder HA558 (Sum[330],Sum[331],Sum[557],Carry_out[557]);
  FullAdder FA559 (Sum[21],Carry_out[330],Carry_out[331],Sum[558],Carry_out[558]);
  HalfAdder HA560 (Sum[332],Sum[333],Sum[559],Carry_out[559]);
  FullAdder FA561 (Carry_out[332],Carry_out[333],Sum[334],Sum[560],Carry_out[560]);
  HalfAdder HA562 (Sum[335],Sum[336],Sum[561],Carry_out[561]);
  FullAdder FA563 (Carry_out[334],Carry_out[335],Carry_out[336],Sum[562],Carry_out[562]);
  FullAdder FA564 (Sum[337],Sum[338],Sum[339],Sum[563],Carry_out[563]);
  FullAdder FA565 (Carry_out[337],Carry_out[338],Carry_out[339],Sum[564],Carry_out[564]);
  FullAdder FA566 (Sum[340],Sum[341],Sum[342],Sum[565],Carry_out[565]);
  FullAdder FA567 (Sum[39],Carry_out[340],Carry_out[341],Sum[566],Carry_out[566]);
  FullAdder FA568 (Carry_out[342],Sum[343],Sum[344],Sum[567],Carry_out[567]);
  FullAdder FA569 (Carry_out[343],Carry_out[344],Carry_out[345],Sum[568],Carry_out[568]);
  FullAdder FA570 (Sum[346],Sum[347],Sum[348],Sum[569],Carry_out[569]);
  FullAdder FA571 (Carry_out[346],Carry_out[347],Carry_out[348],Sum[570],Carry_out[570]);
  FullAdder FA572 (Carry_out[349],Sum[350],Sum[351],Sum[571],Carry_out[571]);
  HalfAdder HA573 (Sum[352],Sum[353],Sum[572],Carry_out[572]);
  FullAdder FA574 (Carry_out[350],Carry_out[351],Carry_out[352],Sum[573],Carry_out[573]);
  FullAdder FA575 (Carry_out[353],Sum[354],Sum[355],Sum[574],Carry_out[574]);
  HalfAdder HA576 (Sum[356],Sum[357],Sum[575],Carry_out[575]);
  FullAdder FA577 (Sum[62],Carry_out[354],Carry_out[355],Sum[576],Carry_out[576]);
  FullAdder FA578 (Carry_out[356],Carry_out[357],Sum[358],Sum[577],Carry_out[577]);
  FullAdder FA579 (Sum[359],Sum[360],Sum[361],Sum[578],Carry_out[578]);
  FullAdder FA580 (Sum[69],Carry_out[358],Carry_out[359],Sum[579],Carry_out[579]);
  FullAdder FA581 (Carry_out[360],Carry_out[361],Sum[362],Sum[580],Carry_out[580]);
  FullAdder FA582 (Sum[363],Sum[364],Sum[365],Sum[581],Carry_out[581]);
  FullAdder FA583 (Carry_out[362],Carry_out[363],Carry_out[364],Sum[582],Carry_out[582]);
  FullAdder FA584 (Carry_out[365],Sum[366],Sum[367],Sum[583],Carry_out[583]);
  FullAdder FA585 (Sum[368],Sum[369],Sum[370],Sum[584],Carry_out[584]);
  FullAdder FA586 (Carry_out[366],Carry_out[367],Carry_out[368],Sum[585],Carry_out[585]);
  FullAdder FA587 (Carry_out[369],Carry_out[370],Sum[371],Sum[586],Carry_out[586]);
  FullAdder FA588 (Sum[372],Sum[373],Sum[374],Sum[587],Carry_out[587]);
  FullAdder FA589 (Carry_out[371],Carry_out[372],Carry_out[373],Sum[588],Carry_out[588]);
  FullAdder FA590 (Carry_out[374],Carry_out[375],Sum[376],Sum[589],Carry_out[589]);
  FullAdder FA591 (Sum[377],Sum[378],Sum[379],Sum[590],Carry_out[590]);
  FullAdder FA592 (Sum[99],Carry_out[376],Carry_out[377],Sum[591],Carry_out[591]);
  FullAdder FA593 (Carry_out[378],Carry_out[379],Carry_out[380],Sum[592],Carry_out[592]);
  FullAdder FA594 (Sum[381],Sum[382],Sum[383],Sum[593],Carry_out[593]);
  HalfAdder HA595 (Sum[384],Sum[385],Sum[594],Carry_out[594]);
  FullAdder FA596 (Carry_out[381],Carry_out[382],Carry_out[383],Sum[595],Carry_out[595]);
  FullAdder FA597 (Carry_out[384],Carry_out[385],Sum[386],Sum[596],Carry_out[596]);
  FullAdder FA598 (Sum[387],Sum[388],Sum[389],Sum[597],Carry_out[597]);
  HalfAdder HA599 (Sum[390],Sum[391],Sum[598],Carry_out[598]);
  FullAdder FA600 (Carry_out[386],Carry_out[387],Carry_out[388],Sum[599],Carry_out[599]);
  FullAdder FA601 (Carry_out[389],Carry_out[390],Carry_out[391],Sum[600],Carry_out[600]);
  FullAdder FA602 (Sum[392],Sum[393],Sum[394],Sum[601],Carry_out[601]);
  FullAdder FA603 (Sum[395],Sum[396],Sum[397],Sum[602],Carry_out[602]);
  FullAdder FA604 (Carry_out[392],Carry_out[393],Carry_out[394],Sum[603],Carry_out[603]);
  FullAdder FA605 (Carry_out[395],Carry_out[396],Carry_out[397],Sum[604],Carry_out[604]);
  FullAdder FA606 (Sum[398],Sum[399],Sum[400],Sum[605],Carry_out[605]);
  FullAdder FA607 (Sum[401],Sum[402],Sum[403],Sum[606],Carry_out[606]);
  FullAdder FA608 (Sum[134],Carry_out[398],Carry_out[399],Sum[607],Carry_out[607]);
  FullAdder FA609 (Carry_out[400],Carry_out[401],Carry_out[402],Sum[608],Carry_out[608]);
  FullAdder FA610 (Carry_out[403],Sum[404],Sum[405],Sum[609],Carry_out[609]);
  FullAdder FA611 (Sum[406],Sum[407],Sum[408],Sum[610],Carry_out[610]);
  FullAdder FA612 (Sum[144],Carry_out[404],Carry_out[405],Sum[611],Carry_out[611]);
  FullAdder FA613 (Carry_out[406],Carry_out[407],Carry_out[408],Sum[612],Carry_out[612]);
  FullAdder FA614 (Carry_out[409],Sum[410],Sum[411],Sum[613],Carry_out[613]);
  FullAdder FA615 (Sum[412],Sum[413],Sum[414],Sum[614],Carry_out[614]);
  FullAdder FA616 (Carry_out[410],Carry_out[411],Carry_out[412],Sum[615],Carry_out[615]);
  FullAdder FA617 (Carry_out[413],Carry_out[414],Carry_out[415],Sum[616],Carry_out[616]);
  FullAdder FA618 (Sum[416],Sum[417],Sum[418],Sum[617],Carry_out[617]);
  FullAdder FA619 (Sum[419],Sum[420],Sum[421],Sum[618],Carry_out[618]);
  FullAdder FA620 (Carry_out[416],Carry_out[417],Carry_out[418],Sum[619],Carry_out[619]);
  FullAdder FA621 (Carry_out[419],Carry_out[420],Carry_out[421],Sum[620],Carry_out[620]);
  FullAdder FA622 (Carry_out[422],Sum[423],Sum[424],Sum[621],Carry_out[621]);
  FullAdder FA623 (Sum[425],Sum[426],Sum[427],Sum[622],Carry_out[622]);
  HalfAdder HA624 (Sum[428],Sum[429],Sum[623],Carry_out[623]);
  FullAdder FA625 (Sum[174],Carry_out[423],Carry_out[424],Sum[624],Carry_out[624]);
  FullAdder FA626 (Carry_out[425],Carry_out[426],Carry_out[427],Sum[625],Carry_out[625]);
  FullAdder FA627 (Carry_out[428],Carry_out[429],Sum[430],Sum[626],Carry_out[626]);
  FullAdder FA628 (Sum[431],Sum[432],Sum[433],Sum[627],Carry_out[627]);
  FullAdder FA629 (Sum[434],Sum[435],Sum[436],Sum[628],Carry_out[628]);
  FullAdder FA630 (Sum[184],Carry_out[430],Carry_out[431],Sum[629],Carry_out[629]);
  FullAdder FA631 (Carry_out[432],Carry_out[433],Carry_out[434],Sum[630],Carry_out[630]);
  FullAdder FA632 (Carry_out[435],Carry_out[436],Sum[437],Sum[631],Carry_out[631]);
  FullAdder FA633 (Sum[438],Sum[439],Sum[440],Sum[632],Carry_out[632]);
  FullAdder FA634 (Sum[441],Sum[442],Sum[443],Sum[633],Carry_out[633]);
  FullAdder FA635 (Sum[193],Carry_out[437],Carry_out[438],Sum[634],Carry_out[634]);
  FullAdder FA636 (Carry_out[439],Carry_out[440],Carry_out[441],Sum[635],Carry_out[635]);
  FullAdder FA637 (Carry_out[442],Carry_out[443],Sum[444],Sum[636],Carry_out[636]);
  FullAdder FA638 (Sum[445],Sum[446],Sum[447],Sum[637],Carry_out[637]);
  FullAdder FA639 (Sum[448],Sum[449],Sum[450],Sum[638],Carry_out[638]);
  FullAdder FA640 (Sum[201],Sum[202],Carry_out[444],Sum[639],Carry_out[639]);
  FullAdder FA641 (Carry_out[445],Carry_out[446],Carry_out[447],Sum[640],Carry_out[640]);
  FullAdder FA642 (Carry_out[448],Carry_out[449],Carry_out[450],Sum[641],Carry_out[641]);
  FullAdder FA643 (Sum[451],Sum[452],Sum[453],Sum[642],Carry_out[642]);
  FullAdder FA644 (Sum[454],Sum[455],Sum[456],Sum[643],Carry_out[643]);
  FullAdder FA645 (Sum[210],Sum[211],Carry_out[451],Sum[644],Carry_out[644]);
  FullAdder FA646 (Carry_out[452],Carry_out[453],Carry_out[454],Sum[645],Carry_out[645]);
  FullAdder FA647 (Carry_out[455],Carry_out[456],Sum[457],Sum[646],Carry_out[646]);
  FullAdder FA648 (Sum[458],Sum[459],Sum[460],Sum[647],Carry_out[647]);
  HalfAdder HA649 (Sum[461],Sum[462],Sum[648],Carry_out[648]);
  FullAdder FA650 (Sum[218],Sum[219],Carry_out[457],Sum[649],Carry_out[649]);
  FullAdder FA651 (Carry_out[458],Carry_out[459],Carry_out[460],Sum[650],Carry_out[650]);
  FullAdder FA652 (Carry_out[461],Carry_out[462],Sum[463],Sum[651],Carry_out[651]);
  FullAdder FA653 (Sum[464],Sum[465],Sum[466],Sum[652],Carry_out[652]);
  HalfAdder HA654 (Sum[467],Sum[468],Sum[653],Carry_out[653]);
  FullAdder FA655 (Sum[227],Carry_out[463],Carry_out[464],Sum[654],Carry_out[654]);
  FullAdder FA656 (Carry_out[465],Carry_out[466],Carry_out[467],Sum[655],Carry_out[655]);
  FullAdder FA657 (Carry_out[468],Sum[469],Sum[470],Sum[656],Carry_out[656]);
  FullAdder FA658 (Sum[471],Sum[472],Sum[473],Sum[657],Carry_out[657]);
  FullAdder FA659 (Sum[235],Carry_out[469],Carry_out[470],Sum[658],Carry_out[658]);
  FullAdder FA660 (Carry_out[471],Carry_out[472],Carry_out[473],Sum[659],Carry_out[659]);
  FullAdder FA661 (Carry_out[474],Sum[475],Sum[476],Sum[660],Carry_out[660]);
  FullAdder FA662 (Sum[477],Sum[478],Sum[479],Sum[661],Carry_out[661]);
  FullAdder FA663 (Sum[242],Carry_out[475],Carry_out[476],Sum[662],Carry_out[662]);
  FullAdder FA664 (Carry_out[477],Carry_out[478],Carry_out[479],Sum[663],Carry_out[663]);
  FullAdder FA665 (Carry_out[480],Sum[481],Sum[482],Sum[664],Carry_out[664]);
  FullAdder FA666 (Sum[483],Sum[484],Sum[485],Sum[665],Carry_out[665]);
  FullAdder FA667 (Sum[249],Carry_out[481],Carry_out[482],Sum[666],Carry_out[666]);
  FullAdder FA668 (Carry_out[483],Carry_out[484],Carry_out[485],Sum[667],Carry_out[667]);
  FullAdder FA669 (Carry_out[486],Sum[487],Sum[488],Sum[668],Carry_out[668]);
  FullAdder FA670 (Sum[489],Sum[490],Sum[491],Sum[669],Carry_out[669]);
  FullAdder FA671 (Sum[256],Carry_out[487],Carry_out[488],Sum[670],Carry_out[670]);
  FullAdder FA672 (Carry_out[489],Carry_out[490],Carry_out[491],Sum[671],Carry_out[671]);
  FullAdder FA673 (Sum[492],Sum[493],Sum[494],Sum[672],Carry_out[672]);
  HalfAdder HA674 (Sum[495],Sum[496],Sum[673],Carry_out[673]);
  FullAdder FA675 (Sum[262],Carry_out[492],Carry_out[493],Sum[674],Carry_out[674]);
  FullAdder FA676 (Carry_out[494],Carry_out[495],Carry_out[496],Sum[675],Carry_out[675]);
  FullAdder FA677 (Sum[497],Sum[498],Sum[499],Sum[676],Carry_out[676]);
  HalfAdder HA678 (Sum[500],Sum[501],Sum[677],Carry_out[677]);
  FullAdder FA679 (Sum[267],Sum[268],Carry_out[497],Sum[678],Carry_out[678]);
  FullAdder FA680 (Carry_out[498],Carry_out[499],Carry_out[500],Sum[679],Carry_out[679]);
  FullAdder FA681 (Carry_out[501],Sum[502],Sum[503],Sum[680],Carry_out[680]);
  HalfAdder HA682 (Sum[504],Sum[505],Sum[681],Carry_out[681]);
  FullAdder FA683 (Sum[273],Sum[274],Carry_out[502],Sum[682],Carry_out[682]);
  FullAdder FA684 (Carry_out[503],Carry_out[504],Carry_out[505],Sum[683],Carry_out[683]);
  FullAdder FA685 (Sum[506],Sum[507],Sum[508],Sum[684],Carry_out[684]);
  FullAdder FA686 (Sum[278],Sum[279],Carry_out[506],Sum[685],Carry_out[685]);
  FullAdder FA687 (Carry_out[507],Carry_out[508],Carry_out[509],Sum[686],Carry_out[686]);
  FullAdder FA688 (Sum[510],Sum[511],Sum[512],Sum[687],Carry_out[687]);
  FullAdder FA689 (Sum[284],Carry_out[510],Carry_out[511],Sum[688],Carry_out[688]);
  FullAdder FA690 (Carry_out[512],Carry_out[513],Sum[514],Sum[689],Carry_out[689]);
  FullAdder FA691 (Sum[515],Sum[516],Sum[517],Sum[690],Carry_out[690]);
  FullAdder FA692 (Sum[289],Carry_out[514],Carry_out[515],Sum[691],Carry_out[691]);
  FullAdder FA693 (Carry_out[516],Carry_out[517],Sum[518],Sum[692],Carry_out[692]);
  FullAdder FA694 (Sum[519],Sum[520],Sum[521],Sum[693],Carry_out[693]);
  FullAdder FA695 (Sum[293],Carry_out[518],Carry_out[519],Sum[694],Carry_out[694]);
  FullAdder FA696 (Carry_out[520],Carry_out[521],Sum[522],Sum[695],Carry_out[695]);
  FullAdder FA697 (Sum[523],Sum[524],Sum[525],Sum[696],Carry_out[696]);
  FullAdder FA698 (Sum[297],Carry_out[522],Carry_out[523],Sum[697],Carry_out[697]);
  FullAdder FA699 (Carry_out[524],Carry_out[525],Sum[526],Sum[698],Carry_out[698]);
  HalfAdder HA700 (Sum[527],Sum[528],Sum[699],Carry_out[699]);
  FullAdder FA701 (Sum[301],Carry_out[526],Carry_out[527],Sum[700],Carry_out[700]);
  FullAdder FA702 (Carry_out[528],Sum[529],Sum[530],Sum[701],Carry_out[701]);
  FullAdder FA703 (Sum[304],Carry_out[529],Carry_out[530],Sum[702],Carry_out[702]);
  FullAdder FA704 (Carry_out[531],Sum[532],Sum[533],Sum[703],Carry_out[703]);
  FullAdder FA705 (Sum[306],Sum[307],Carry_out[532],Sum[704],Carry_out[704]);
  FullAdder FA706 (Carry_out[533],Carry_out[534],Sum[535],Sum[705],Carry_out[705]);
  FullAdder FA707 (Sum[309],Sum[310],Carry_out[535],Sum[706],Carry_out[706]);
  FullAdder FA708 (Carry_out[536],Sum[537],Sum[538],Sum[707],Carry_out[707]);
  FullAdder FA709 (Sum[311],Sum[312],Carry_out[537],Sum[708],Carry_out[708]);
  FullAdder FA710 (Carry_out[538],Sum[539],Sum[540],Sum[709],Carry_out[709]);
  FullAdder FA711 (Sum[314],Carry_out[539],Carry_out[540],Sum[710],Carry_out[710]);
  HalfAdder HA712 (Sum[541],Sum[542],Sum[711],Carry_out[711]);
  FullAdder FA713 (Sum[316],Carry_out[541],Carry_out[542],Sum[712],Carry_out[712]);
  HalfAdder HA714 (Sum[543],Sum[544],Sum[713],Carry_out[713]);
  FullAdder FA715 (Sum[317],Carry_out[543],Carry_out[544],Sum[714],Carry_out[714]);
  HalfAdder HA716 (Sum[545],Sum[546],Sum[715],Carry_out[715]);
  FullAdder FA717 (Sum[318],Carry_out[545],Carry_out[546],Sum[716],Carry_out[716]);
  FullAdder FA718 (Sum[319],Carry_out[547],Sum[548],Sum[717],Carry_out[717]);
  FullAdder FA719 (Carry_out[319],Carry_out[548],Sum[549],Sum[718],Carry_out[718]);
  FullAdder FA720 (Partial_Product[30][31],Partial_Product[31][30],Carry_out[549],Sum[719],Carry_out[719]);
  HalfAdder HA721 (Carry_out[550],Sum[551],Sum[720],Carry_out[720]);
  HalfAdder HA722 (Carry_out[551],Sum[552],Sum[721],Carry_out[721]);
  HalfAdder HA723 (Carry_out[552],Sum[553],Sum[722],Carry_out[722]);
  FullAdder FA724 (Sum[327],Carry_out[553],Sum[554],Sum[723],Carry_out[723]);
  FullAdder FA725 (Sum[329],Carry_out[554],Sum[555],Sum[724],Carry_out[724]);
  FullAdder FA726 (Carry_out[555],Sum[556],Sum[557],Sum[725],Carry_out[725]);
  FullAdder FA727 (Carry_out[556],Carry_out[557],Sum[558],Sum[726],Carry_out[726]);
  FullAdder FA728 (Carry_out[558],Carry_out[559],Sum[560],Sum[727],Carry_out[727]);
  FullAdder FA729 (Carry_out[560],Carry_out[561],Sum[562],Sum[728],Carry_out[728]);
  FullAdder FA730 (Carry_out[562],Carry_out[563],Sum[564],Sum[729],Carry_out[729]);
  FullAdder FA731 (Sum[345],Carry_out[564],Carry_out[565],Sum[730],Carry_out[730]);
  HalfAdder HA732 (Sum[566],Sum[567],Sum[731],Carry_out[731]);
  FullAdder FA733 (Sum[349],Carry_out[566],Carry_out[567],Sum[732],Carry_out[732]);
  HalfAdder HA734 (Sum[568],Sum[569],Sum[733],Carry_out[733]);
  FullAdder FA735 (Carry_out[568],Carry_out[569],Sum[570],Sum[734],Carry_out[734]);
  HalfAdder HA736 (Sum[571],Sum[572],Sum[735],Carry_out[735]);
  FullAdder FA737 (Carry_out[570],Carry_out[571],Carry_out[572],Sum[736],Carry_out[736]);
  FullAdder FA738 (Sum[573],Sum[574],Sum[575],Sum[737],Carry_out[737]);
  FullAdder FA739 (Carry_out[573],Carry_out[574],Carry_out[575],Sum[738],Carry_out[738]);
  FullAdder FA740 (Sum[576],Sum[577],Sum[578],Sum[739],Carry_out[739]);
  FullAdder FA741 (Carry_out[576],Carry_out[577],Carry_out[578],Sum[740],Carry_out[740]);
  FullAdder FA742 (Sum[579],Sum[580],Sum[581],Sum[741],Carry_out[741]);
  FullAdder FA743 (Carry_out[579],Carry_out[580],Carry_out[581],Sum[742],Carry_out[742]);
  FullAdder FA744 (Sum[582],Sum[583],Sum[584],Sum[743],Carry_out[743]);
  FullAdder FA745 (Sum[375],Carry_out[582],Carry_out[583],Sum[744],Carry_out[744]);
  FullAdder FA746 (Carry_out[584],Sum[585],Sum[586],Sum[745],Carry_out[745]);
  FullAdder FA747 (Sum[380],Carry_out[585],Carry_out[586],Sum[746],Carry_out[746]);
  FullAdder FA748 (Carry_out[587],Sum[588],Sum[589],Sum[747],Carry_out[747]);
  FullAdder FA749 (Carry_out[588],Carry_out[589],Carry_out[590],Sum[748],Carry_out[748]);
  FullAdder FA750 (Sum[591],Sum[592],Sum[593],Sum[749],Carry_out[749]);
  FullAdder FA751 (Carry_out[591],Carry_out[592],Carry_out[593],Sum[750],Carry_out[750]);
  FullAdder FA752 (Carry_out[594],Sum[595],Sum[596],Sum[751],Carry_out[751]);
  HalfAdder HA753 (Sum[597],Sum[598],Sum[752],Carry_out[752]);
  FullAdder FA754 (Carry_out[595],Carry_out[596],Carry_out[597],Sum[753],Carry_out[753]);
  FullAdder FA755 (Carry_out[598],Sum[599],Sum[600],Sum[754],Carry_out[754]);
  HalfAdder HA756 (Sum[601],Sum[602],Sum[755],Carry_out[755]);
  FullAdder FA757 (Carry_out[599],Carry_out[600],Carry_out[601],Sum[756],Carry_out[756]);
  FullAdder FA758 (Carry_out[602],Sum[603],Sum[604],Sum[757],Carry_out[757]);
  HalfAdder HA759 (Sum[605],Sum[606],Sum[758],Carry_out[758]);
  FullAdder FA760 (Sum[409],Carry_out[603],Carry_out[604],Sum[759],Carry_out[759]);
  FullAdder FA761 (Carry_out[605],Carry_out[606],Sum[607],Sum[760],Carry_out[760]);
  FullAdder FA762 (Sum[608],Sum[609],Sum[610],Sum[761],Carry_out[761]);
  FullAdder FA763 (Sum[415],Carry_out[607],Carry_out[608],Sum[762],Carry_out[762]);
  FullAdder FA764 (Carry_out[609],Carry_out[610],Sum[611],Sum[763],Carry_out[763]);
  FullAdder FA765 (Sum[612],Sum[613],Sum[614],Sum[764],Carry_out[764]);
  FullAdder FA766 (Sum[422],Carry_out[611],Carry_out[612],Sum[765],Carry_out[765]);
  FullAdder FA767 (Carry_out[613],Carry_out[614],Sum[615],Sum[766],Carry_out[766]);
  FullAdder FA768 (Sum[616],Sum[617],Sum[618],Sum[767],Carry_out[767]);
  FullAdder FA769 (Carry_out[615],Carry_out[616],Carry_out[617],Sum[768],Carry_out[768]);
  FullAdder FA770 (Carry_out[618],Sum[619],Sum[620],Sum[769],Carry_out[769]);
  FullAdder FA771 (Sum[621],Sum[622],Sum[623],Sum[770],Carry_out[770]);
  FullAdder FA772 (Carry_out[619],Carry_out[620],Carry_out[621],Sum[771],Carry_out[771]);
  FullAdder FA773 (Carry_out[622],Carry_out[623],Sum[624],Sum[772],Carry_out[772]);
  FullAdder FA774 (Sum[625],Sum[626],Sum[627],Sum[773],Carry_out[773]);
  FullAdder FA775 (Carry_out[624],Carry_out[625],Carry_out[626],Sum[774],Carry_out[774]);
  FullAdder FA776 (Carry_out[627],Carry_out[628],Sum[629],Sum[775],Carry_out[775]);
  FullAdder FA777 (Sum[630],Sum[631],Sum[632],Sum[776],Carry_out[776]);
  FullAdder FA778 (Carry_out[629],Carry_out[630],Carry_out[631],Sum[777],Carry_out[777]);
  FullAdder FA779 (Carry_out[632],Carry_out[633],Sum[634],Sum[778],Carry_out[778]);
  FullAdder FA780 (Sum[635],Sum[636],Sum[637],Sum[779],Carry_out[779]);
  FullAdder FA781 (Carry_out[634],Carry_out[635],Carry_out[636],Sum[780],Carry_out[780]);
  FullAdder FA782 (Carry_out[637],Carry_out[638],Sum[639],Sum[781],Carry_out[781]);
  FullAdder FA783 (Sum[640],Sum[641],Sum[642],Sum[782],Carry_out[782]);
  FullAdder FA784 (Carry_out[639],Carry_out[640],Carry_out[641],Sum[783],Carry_out[783]);
  FullAdder FA785 (Carry_out[642],Carry_out[643],Sum[644],Sum[784],Carry_out[784]);
  FullAdder FA786 (Sum[645],Sum[646],Sum[647],Sum[785],Carry_out[785]);
  FullAdder FA787 (Carry_out[644],Carry_out[645],Carry_out[646],Sum[786],Carry_out[786]);
  FullAdder FA788 (Carry_out[647],Carry_out[648],Sum[649],Sum[787],Carry_out[787]);
  FullAdder FA789 (Sum[650],Sum[651],Sum[652],Sum[788],Carry_out[788]);
  FullAdder FA790 (Sum[474],Carry_out[649],Carry_out[650],Sum[789],Carry_out[789]);
  FullAdder FA791 (Carry_out[651],Carry_out[652],Carry_out[653],Sum[790],Carry_out[790]);
  FullAdder FA792 (Sum[654],Sum[655],Sum[656],Sum[791],Carry_out[791]);
  FullAdder FA793 (Sum[480],Carry_out[654],Carry_out[655],Sum[792],Carry_out[792]);
  FullAdder FA794 (Carry_out[656],Carry_out[657],Sum[658],Sum[793],Carry_out[793]);
  HalfAdder HA795 (Sum[659],Sum[660],Sum[794],Carry_out[794]);
  FullAdder FA796 (Sum[486],Carry_out[658],Carry_out[659],Sum[795],Carry_out[795]);
  FullAdder FA797 (Carry_out[660],Carry_out[661],Sum[662],Sum[796],Carry_out[796]);
  HalfAdder HA798 (Sum[663],Sum[664],Sum[797],Carry_out[797]);
  FullAdder FA799 (Carry_out[662],Carry_out[663],Carry_out[664],Sum[798],Carry_out[798]);
  FullAdder FA800 (Carry_out[665],Sum[666],Sum[667],Sum[799],Carry_out[799]);
  FullAdder FA801 (Carry_out[666],Carry_out[667],Carry_out[668],Sum[800],Carry_out[800]);
  FullAdder FA802 (Carry_out[669],Sum[670],Sum[671],Sum[801],Carry_out[801]);
  FullAdder FA803 (Carry_out[670],Carry_out[671],Carry_out[672],Sum[802],Carry_out[802]);
  FullAdder FA804 (Carry_out[673],Sum[674],Sum[675],Sum[803],Carry_out[803]);
  FullAdder FA805 (Carry_out[674],Carry_out[675],Carry_out[676],Sum[804],Carry_out[804]);
  FullAdder FA806 (Carry_out[677],Sum[678],Sum[679],Sum[805],Carry_out[805]);
  FullAdder FA807 (Sum[509],Carry_out[678],Carry_out[679],Sum[806],Carry_out[806]);
  FullAdder FA808 (Carry_out[680],Carry_out[681],Sum[682],Sum[807],Carry_out[807]);
  FullAdder FA809 (Sum[513],Carry_out[682],Carry_out[683],Sum[808],Carry_out[808]);
  FullAdder FA810 (Carry_out[684],Sum[685],Sum[686],Sum[809],Carry_out[809]);
  FullAdder FA811 (Carry_out[685],Carry_out[686],Carry_out[687],Sum[810],Carry_out[810]);
  HalfAdder HA812 (Sum[688],Sum[689],Sum[811],Carry_out[811]);
  FullAdder FA813 (Carry_out[688],Carry_out[689],Carry_out[690],Sum[812],Carry_out[812]);
  HalfAdder HA814 (Sum[691],Sum[692],Sum[813],Carry_out[813]);
  FullAdder FA815 (Carry_out[691],Carry_out[692],Carry_out[693],Sum[814],Carry_out[814]);
  HalfAdder HA816 (Sum[694],Sum[695],Sum[815],Carry_out[815]);
  FullAdder FA817 (Carry_out[694],Carry_out[695],Carry_out[696],Sum[816],Carry_out[816]);
  HalfAdder HA818 (Sum[697],Sum[698],Sum[817],Carry_out[817]);
  FullAdder FA819 (Sum[531],Carry_out[697],Carry_out[698],Sum[818],Carry_out[818]);
  HalfAdder HA820 (Carry_out[699],Sum[700],Sum[819],Carry_out[819]);
  FullAdder FA821 (Sum[534],Carry_out[700],Carry_out[701],Sum[820],Carry_out[820]);
  FullAdder FA822 (Sum[536],Carry_out[702],Carry_out[703],Sum[821],Carry_out[821]);
  FullAdder FA823 (Carry_out[704],Carry_out[705],Sum[706],Sum[822],Carry_out[822]);
  FullAdder FA824 (Carry_out[706],Carry_out[707],Sum[708],Sum[823],Carry_out[823]);
  FullAdder FA825 (Carry_out[708],Carry_out[709],Sum[710],Sum[824],Carry_out[824]);
  FullAdder FA826 (Carry_out[710],Carry_out[711],Sum[712],Sum[825],Carry_out[825]);
  FullAdder FA827 (Carry_out[712],Carry_out[713],Sum[714],Sum[826],Carry_out[826]);
  FullAdder FA828 (Sum[547],Carry_out[714],Carry_out[715],Sum[827],Carry_out[827]);
  HalfAdder HA829 (Carry_out[720],Sum[721],Sum[828],Carry_out[828]);
  HalfAdder HA830 (Carry_out[721],Sum[722],Sum[829],Carry_out[829]);
  HalfAdder HA831 (Carry_out[722],Sum[723],Sum[830],Carry_out[830]);
  HalfAdder HA832 (Carry_out[723],Sum[724],Sum[831],Carry_out[831]);
  HalfAdder HA833 (Carry_out[724],Sum[725],Sum[832],Carry_out[832]);
  FullAdder FA834 (Sum[559],Carry_out[725],Sum[726],Sum[833],Carry_out[833]);
  FullAdder FA835 (Sum[561],Carry_out[726],Sum[727],Sum[834],Carry_out[834]);
  FullAdder FA836 (Sum[563],Carry_out[727],Sum[728],Sum[835],Carry_out[835]);
  FullAdder FA837 (Sum[565],Carry_out[728],Sum[729],Sum[836],Carry_out[836]);
  FullAdder FA838 (Carry_out[729],Sum[730],Sum[731],Sum[837],Carry_out[837]);
  FullAdder FA839 (Carry_out[730],Carry_out[731],Sum[732],Sum[838],Carry_out[838]);
  FullAdder FA840 (Carry_out[732],Carry_out[733],Sum[734],Sum[839],Carry_out[839]);
  FullAdder FA841 (Carry_out[734],Carry_out[735],Sum[736],Sum[840],Carry_out[840]);
  FullAdder FA842 (Carry_out[736],Carry_out[737],Sum[738],Sum[841],Carry_out[841]);
  FullAdder FA843 (Carry_out[738],Carry_out[739],Sum[740],Sum[842],Carry_out[842]);
  FullAdder FA844 (Carry_out[740],Carry_out[741],Sum[742],Sum[843],Carry_out[843]);
  FullAdder FA845 (Sum[587],Carry_out[742],Carry_out[743],Sum[844],Carry_out[844]);
  HalfAdder HA846 (Sum[744],Sum[745],Sum[845],Carry_out[845]);
  FullAdder FA847 (Sum[590],Carry_out[744],Carry_out[745],Sum[846],Carry_out[846]);
  HalfAdder HA848 (Sum[746],Sum[747],Sum[847],Carry_out[847]);
  FullAdder FA849 (Sum[594],Carry_out[746],Carry_out[747],Sum[848],Carry_out[848]);
  HalfAdder HA850 (Sum[748],Sum[749],Sum[849],Carry_out[849]);
  FullAdder FA851 (Carry_out[748],Carry_out[749],Sum[750],Sum[850],Carry_out[850]);
  HalfAdder HA852 (Sum[751],Sum[752],Sum[851],Carry_out[851]);
  FullAdder FA853 (Carry_out[750],Carry_out[751],Carry_out[752],Sum[852],Carry_out[852]);
  FullAdder FA854 (Sum[753],Sum[754],Sum[755],Sum[853],Carry_out[853]);
  FullAdder FA855 (Carry_out[753],Carry_out[754],Carry_out[755],Sum[854],Carry_out[854]);
  FullAdder FA856 (Sum[756],Sum[757],Sum[758],Sum[855],Carry_out[855]);
  FullAdder FA857 (Carry_out[756],Carry_out[757],Carry_out[758],Sum[856],Carry_out[856]);
  FullAdder FA858 (Sum[759],Sum[760],Sum[761],Sum[857],Carry_out[857]);
  FullAdder FA859 (Carry_out[759],Carry_out[760],Carry_out[761],Sum[858],Carry_out[858]);
  FullAdder FA860 (Sum[762],Sum[763],Sum[764],Sum[859],Carry_out[859]);
  FullAdder FA861 (Carry_out[762],Carry_out[763],Carry_out[764],Sum[860],Carry_out[860]);
  FullAdder FA862 (Sum[765],Sum[766],Sum[767],Sum[861],Carry_out[861]);
  FullAdder FA863 (Carry_out[765],Carry_out[766],Carry_out[767],Sum[862],Carry_out[862]);
  FullAdder FA864 (Sum[768],Sum[769],Sum[770],Sum[863],Carry_out[863]);
  FullAdder FA865 (Sum[628],Carry_out[768],Carry_out[769],Sum[864],Carry_out[864]);
  FullAdder FA866 (Carry_out[770],Sum[771],Sum[772],Sum[865],Carry_out[865]);
  FullAdder FA867 (Sum[633],Carry_out[771],Carry_out[772],Sum[866],Carry_out[866]);
  FullAdder FA868 (Carry_out[773],Sum[774],Sum[775],Sum[867],Carry_out[867]);
  FullAdder FA869 (Sum[638],Carry_out[774],Carry_out[775],Sum[868],Carry_out[868]);
  FullAdder FA870 (Carry_out[776],Sum[777],Sum[778],Sum[869],Carry_out[869]);
  FullAdder FA871 (Sum[643],Carry_out[777],Carry_out[778],Sum[870],Carry_out[870]);
  FullAdder FA872 (Carry_out[779],Sum[780],Sum[781],Sum[871],Carry_out[871]);
  FullAdder FA873 (Sum[648],Carry_out[780],Carry_out[781],Sum[872],Carry_out[872]);
  FullAdder FA874 (Carry_out[782],Sum[783],Sum[784],Sum[873],Carry_out[873]);
  FullAdder FA875 (Sum[653],Carry_out[783],Carry_out[784],Sum[874],Carry_out[874]);
  FullAdder FA876 (Carry_out[785],Sum[786],Sum[787],Sum[875],Carry_out[875]);
  FullAdder FA877 (Sum[657],Carry_out[786],Carry_out[787],Sum[876],Carry_out[876]);
  FullAdder FA878 (Carry_out[788],Sum[789],Sum[790],Sum[877],Carry_out[877]);
  FullAdder FA879 (Sum[661],Carry_out[789],Carry_out[790],Sum[878],Carry_out[878]);
  FullAdder FA880 (Carry_out[791],Sum[792],Sum[793],Sum[879],Carry_out[879]);
  FullAdder FA881 (Sum[665],Carry_out[792],Carry_out[793],Sum[880],Carry_out[880]);
  FullAdder FA882 (Carry_out[794],Sum[795],Sum[796],Sum[881],Carry_out[881]);
  FullAdder FA883 (Sum[668],Sum[669],Carry_out[795],Sum[882],Carry_out[882]);
  FullAdder FA884 (Carry_out[796],Carry_out[797],Sum[798],Sum[883],Carry_out[883]);
  FullAdder FA885 (Sum[672],Sum[673],Carry_out[798],Sum[884],Carry_out[884]);
  HalfAdder HA886 (Carry_out[799],Sum[800],Sum[885],Carry_out[885]);
  FullAdder FA887 (Sum[676],Sum[677],Carry_out[800],Sum[886],Carry_out[886]);
  HalfAdder HA888 (Carry_out[801],Sum[802],Sum[887],Carry_out[887]);
  FullAdder FA889 (Sum[680],Sum[681],Carry_out[802],Sum[888],Carry_out[888]);
  HalfAdder HA890 (Carry_out[803],Sum[804],Sum[889],Carry_out[889]);
  FullAdder FA891 (Sum[683],Sum[684],Carry_out[804],Sum[890],Carry_out[890]);
  HalfAdder HA892 (Carry_out[805],Sum[806],Sum[891],Carry_out[891]);
  FullAdder FA893 (Sum[687],Carry_out[806],Carry_out[807],Sum[892],Carry_out[892]);
  FullAdder FA894 (Sum[690],Carry_out[808],Carry_out[809],Sum[893],Carry_out[893]);
  FullAdder FA895 (Sum[693],Carry_out[810],Carry_out[811],Sum[894],Carry_out[894]);
  FullAdder FA896 (Sum[696],Carry_out[812],Carry_out[813],Sum[895],Carry_out[895]);
  FullAdder FA897 (Sum[699],Carry_out[814],Carry_out[815],Sum[896],Carry_out[896]);
  FullAdder FA898 (Sum[701],Carry_out[816],Carry_out[817],Sum[897],Carry_out[897]);
  FullAdder FA899 (Sum[702],Sum[703],Carry_out[818],Sum[898],Carry_out[898]);
  FullAdder FA900 (Sum[704],Sum[705],Carry_out[820],Sum[899],Carry_out[899]);
  HalfAdder HA901 (Sum[707],Carry_out[821],Sum[900],Carry_out[900]);
  HalfAdder HA902 (Sum[709],Carry_out[822],Sum[901],Carry_out[901]);
  HalfAdder HA903 (Sum[711],Carry_out[823],Sum[902],Carry_out[902]);
  HalfAdder HA904 (Sum[713],Carry_out[824],Sum[903],Carry_out[903]);
  HalfAdder HA905 (Sum[715],Carry_out[825],Sum[904],Carry_out[904]);
  HalfAdder HA906 (Sum[716],Carry_out[826],Sum[905],Carry_out[905]);
  HalfAdder HA907 (Carry_out[716],Sum[717],Sum[906],Carry_out[906]);
  HalfAdder HA908 (Carry_out[828],Sum[829],Sum[907],Carry_out[907]);
  HalfAdder HA909 (Carry_out[829],Sum[830],Sum[908],Carry_out[908]);
  HalfAdder HA910 (Carry_out[830],Sum[831],Sum[909],Carry_out[909]);
  HalfAdder HA911 (Carry_out[831],Sum[832],Sum[910],Carry_out[910]);
  HalfAdder HA912 (Carry_out[832],Sum[833],Sum[911],Carry_out[911]);
  HalfAdder HA913 (Carry_out[833],Sum[834],Sum[912],Carry_out[912]);
  HalfAdder HA914 (Carry_out[834],Sum[835],Sum[913],Carry_out[913]);
  HalfAdder HA915 (Carry_out[835],Sum[836],Sum[914],Carry_out[914]);
  HalfAdder HA916 (Carry_out[836],Sum[837],Sum[915],Carry_out[915]);
  FullAdder FA917 (Sum[733],Carry_out[837],Sum[838],Sum[916],Carry_out[916]);
  FullAdder FA918 (Sum[735],Carry_out[838],Sum[839],Sum[917],Carry_out[917]);
  FullAdder FA919 (Sum[737],Carry_out[839],Sum[840],Sum[918],Carry_out[918]);
  FullAdder FA920 (Sum[739],Carry_out[840],Sum[841],Sum[919],Carry_out[919]);
  FullAdder FA921 (Sum[741],Carry_out[841],Sum[842],Sum[920],Carry_out[920]);
  FullAdder FA922 (Sum[743],Carry_out[842],Sum[843],Sum[921],Carry_out[921]);
  FullAdder FA923 (Carry_out[843],Sum[844],Sum[845],Sum[922],Carry_out[922]);
  FullAdder FA924 (Carry_out[844],Carry_out[845],Sum[846],Sum[923],Carry_out[923]);
  FullAdder FA925 (Carry_out[846],Carry_out[847],Sum[848],Sum[924],Carry_out[924]);
  FullAdder FA926 (Carry_out[848],Carry_out[849],Sum[850],Sum[925],Carry_out[925]);
  FullAdder FA927 (Carry_out[850],Carry_out[851],Sum[852],Sum[926],Carry_out[926]);
  FullAdder FA928 (Carry_out[852],Carry_out[853],Sum[854],Sum[927],Carry_out[927]);
  FullAdder FA929 (Carry_out[854],Carry_out[855],Sum[856],Sum[928],Carry_out[928]);
  FullAdder FA930 (Carry_out[856],Carry_out[857],Sum[858],Sum[929],Carry_out[929]);
  FullAdder FA931 (Carry_out[858],Carry_out[859],Sum[860],Sum[930],Carry_out[930]);
  FullAdder FA932 (Carry_out[860],Carry_out[861],Sum[862],Sum[931],Carry_out[931]);
  FullAdder FA933 (Sum[773],Carry_out[862],Carry_out[863],Sum[932],Carry_out[932]);
  FullAdder FA934 (Sum[776],Carry_out[864],Carry_out[865],Sum[933],Carry_out[933]);
  FullAdder FA935 (Sum[779],Carry_out[866],Carry_out[867],Sum[934],Carry_out[934]);
  FullAdder FA936 (Sum[782],Carry_out[868],Carry_out[869],Sum[935],Carry_out[935]);
  FullAdder FA937 (Sum[785],Carry_out[870],Carry_out[871],Sum[936],Carry_out[936]);
  FullAdder FA938 (Sum[788],Carry_out[872],Carry_out[873],Sum[937],Carry_out[937]);
  FullAdder FA939 (Sum[791],Carry_out[874],Carry_out[875],Sum[938],Carry_out[938]);
  FullAdder FA940 (Sum[794],Carry_out[876],Carry_out[877],Sum[939],Carry_out[939]);
  FullAdder FA941 (Sum[797],Carry_out[878],Carry_out[879],Sum[940],Carry_out[940]);
  FullAdder FA942 (Sum[799],Carry_out[880],Carry_out[881],Sum[941],Carry_out[941]);
  FullAdder FA943 (Sum[801],Carry_out[882],Carry_out[883],Sum[942],Carry_out[942]);
  FullAdder FA944 (Sum[803],Carry_out[884],Carry_out[885],Sum[943],Carry_out[943]);
  FullAdder FA945 (Sum[805],Carry_out[886],Carry_out[887],Sum[944],Carry_out[944]);
  FullAdder FA946 (Sum[807],Carry_out[888],Carry_out[889],Sum[945],Carry_out[945]);
  FullAdder FA947 (Sum[808],Sum[809],Carry_out[890],Sum[946],Carry_out[946]);
  HalfAdder HA948 (Sum[810],Sum[811],Sum[947],Carry_out[947]);
  HalfAdder HA949 (Sum[812],Sum[813],Sum[948],Carry_out[948]);
  HalfAdder HA950 (Sum[814],Sum[815],Sum[949],Carry_out[949]);
  HalfAdder HA951 (Sum[816],Sum[817],Sum[950],Carry_out[950]);
  HalfAdder HA952 (Sum[818],Sum[819],Sum[951],Carry_out[951]);
  HalfAdder HA953 (Carry_out[819],Sum[820],Sum[952],Carry_out[952]);
  HalfAdder HA954 (Carry_out[907],Sum[908],Sum[953],Carry_out[953]);
  HalfAdder HA955 (Carry_out[908],Sum[909],Sum[954],Carry_out[954]);
  HalfAdder HA956 (Carry_out[909],Sum[910],Sum[955],Carry_out[955]);
  HalfAdder HA957 (Carry_out[910],Sum[911],Sum[956],Carry_out[956]);
  HalfAdder HA958 (Carry_out[911],Sum[912],Sum[957],Carry_out[957]);
  HalfAdder HA959 (Carry_out[912],Sum[913],Sum[958],Carry_out[958]);
  HalfAdder HA960 (Carry_out[913],Sum[914],Sum[959],Carry_out[959]);
  HalfAdder HA961 (Carry_out[914],Sum[915],Sum[960],Carry_out[960]);
  HalfAdder HA962 (Carry_out[915],Sum[916],Sum[961],Carry_out[961]);
  HalfAdder HA963 (Carry_out[916],Sum[917],Sum[962],Carry_out[962]);
  HalfAdder HA964 (Carry_out[917],Sum[918],Sum[963],Carry_out[963]);
  HalfAdder HA965 (Carry_out[918],Sum[919],Sum[964],Carry_out[964]);
  HalfAdder HA966 (Carry_out[919],Sum[920],Sum[965],Carry_out[965]);
  HalfAdder HA967 (Carry_out[920],Sum[921],Sum[966],Carry_out[966]);
  HalfAdder HA968 (Carry_out[921],Sum[922],Sum[967],Carry_out[967]);
  FullAdder FA969 (Sum[847],Carry_out[922],Sum[923],Sum[968],Carry_out[968]);
  FullAdder FA970 (Sum[849],Carry_out[923],Sum[924],Sum[969],Carry_out[969]);
  FullAdder FA971 (Sum[851],Carry_out[924],Sum[925],Sum[970],Carry_out[970]);
  FullAdder FA972 (Sum[853],Carry_out[925],Sum[926],Sum[971],Carry_out[971]);
  FullAdder FA973 (Sum[855],Carry_out[926],Sum[927],Sum[972],Carry_out[972]);
  FullAdder FA974 (Sum[857],Carry_out[927],Sum[928],Sum[973],Carry_out[973]);
  FullAdder FA975 (Sum[859],Carry_out[928],Sum[929],Sum[974],Carry_out[974]);
  FullAdder FA976 (Sum[861],Carry_out[929],Sum[930],Sum[975],Carry_out[975]);
  FullAdder FA977 (Sum[863],Carry_out[930],Sum[931],Sum[976],Carry_out[976]);
  FullAdder FA978 (Sum[864],Sum[865],Carry_out[931],Sum[977],Carry_out[977]);
  FullAdder FA979 (Sum[866],Sum[867],Carry_out[932],Sum[978],Carry_out[978]);
  FullAdder FA980 (Sum[868],Sum[869],Carry_out[933],Sum[979],Carry_out[979]);
  FullAdder FA981 (Sum[870],Sum[871],Carry_out[934],Sum[980],Carry_out[980]);
  FullAdder FA982 (Sum[872],Sum[873],Carry_out[935],Sum[981],Carry_out[981]);
  FullAdder FA983 (Sum[874],Sum[875],Carry_out[936],Sum[982],Carry_out[982]);
  FullAdder FA984 (Sum[876],Sum[877],Carry_out[937],Sum[983],Carry_out[983]);
  FullAdder FA985 (Sum[878],Sum[879],Carry_out[938],Sum[984],Carry_out[984]);
  FullAdder FA986 (Sum[880],Sum[881],Carry_out[939],Sum[985],Carry_out[985]);
  FullAdder FA987 (Sum[882],Sum[883],Carry_out[940],Sum[986],Carry_out[986]);
  FullAdder FA988 (Sum[884],Sum[885],Carry_out[941],Sum[987],Carry_out[987]);
  FullAdder FA989 (Sum[886],Sum[887],Carry_out[942],Sum[988],Carry_out[988]);
  FullAdder FA990 (Sum[888],Sum[889],Carry_out[943],Sum[989],Carry_out[989]);
  FullAdder FA991 (Sum[890],Sum[891],Carry_out[944],Sum[990],Carry_out[990]);
  FullAdder FA992 (Carry_out[891],Sum[892],Carry_out[945],Sum[991],Carry_out[991]);
  FullAdder FA993 (Carry_out[892],Sum[893],Carry_out[946],Sum[992],Carry_out[992]);
  FullAdder FA994 (Carry_out[893],Sum[894],Carry_out[947],Sum[993],Carry_out[993]);
  FullAdder FA995 (Carry_out[894],Sum[895],Carry_out[948],Sum[994],Carry_out[994]);
  FullAdder FA996 (Carry_out[895],Sum[896],Carry_out[949],Sum[995],Carry_out[995]);
  FullAdder FA997 (Carry_out[896],Sum[897],Carry_out[950],Sum[996],Carry_out[996]);
  FullAdder FA998 (Carry_out[897],Sum[898],Carry_out[951],Sum[997],Carry_out[997]);
  FullAdder FA999 (Sum[821],Carry_out[898],Sum[899],Sum[998],Carry_out[998]);
  HalfAdder HA1000 (Sum[822],Carry_out[899],Sum[999],Carry_out[999]);
  HalfAdder HA1001 (Sum[823],Carry_out[900],Sum[1000],Carry_out[1000]);
  HalfAdder HA1002 (Sum[824],Carry_out[901],Sum[1001],Carry_out[1001]);
  HalfAdder HA1003 (Sum[825],Carry_out[902],Sum[1002],Carry_out[1002]);
  HalfAdder HA1004 (Sum[826],Carry_out[903],Sum[1003],Carry_out[1003]);
  HalfAdder HA1005 (Sum[827],Carry_out[904],Sum[1004],Carry_out[1004]);
  HalfAdder HA1006 (Carry_out[827],Carry_out[905],Sum[1005],Carry_out[1005]);
  HalfAdder HA1007 (Carry_out[717],Sum[718],Sum[1006],Carry_out[1006]);
  HalfAdder HA1008 (Carry_out[953],Sum[954],Sum[1007],Carry_out[1007]);
  HalfAdder HA1009 (Carry_out[954],Sum[955],Sum[1008],Carry_out[1008]);
  HalfAdder HA1010 (Carry_out[955],Sum[956],Sum[1009],Carry_out[1009]);
  HalfAdder HA1011 (Carry_out[956],Sum[957],Sum[1010],Carry_out[1010]);
  HalfAdder HA1012 (Carry_out[957],Sum[958],Sum[1011],Carry_out[1011]);
  HalfAdder HA1013 (Carry_out[958],Sum[959],Sum[1012],Carry_out[1012]);
  HalfAdder HA1014 (Carry_out[959],Sum[960],Sum[1013],Carry_out[1013]);
  HalfAdder HA1015 (Carry_out[960],Sum[961],Sum[1014],Carry_out[1014]);
  HalfAdder HA1016 (Carry_out[961],Sum[962],Sum[1015],Carry_out[1015]);
  HalfAdder HA1017 (Carry_out[962],Sum[963],Sum[1016],Carry_out[1016]);
  HalfAdder HA1018 (Carry_out[963],Sum[964],Sum[1017],Carry_out[1017]);
  HalfAdder HA1019 (Carry_out[964],Sum[965],Sum[1018],Carry_out[1018]);
  HalfAdder HA1020 (Carry_out[965],Sum[966],Sum[1019],Carry_out[1019]);
  HalfAdder HA1021 (Carry_out[966],Sum[967],Sum[1020],Carry_out[1020]);
  HalfAdder HA1022 (Carry_out[967],Sum[968],Sum[1021],Carry_out[1021]);
  HalfAdder HA1023 (Carry_out[968],Sum[969],Sum[1022],Carry_out[1022]);
  HalfAdder HA1024 (Carry_out[969],Sum[970],Sum[1023],Carry_out[1023]);
  HalfAdder HA1025 (Carry_out[970],Sum[971],Sum[1024],Carry_out[1024]);
  HalfAdder HA1026 (Carry_out[971],Sum[972],Sum[1025],Carry_out[1025]);
  HalfAdder HA1027 (Carry_out[972],Sum[973],Sum[1026],Carry_out[1026]);
  HalfAdder HA1028 (Carry_out[973],Sum[974],Sum[1027],Carry_out[1027]);
  HalfAdder HA1029 (Carry_out[974],Sum[975],Sum[1028],Carry_out[1028]);
  HalfAdder HA1030 (Carry_out[975],Sum[976],Sum[1029],Carry_out[1029]);
  FullAdder FA1031 (Sum[932],Carry_out[976],Sum[977],Sum[1030],Carry_out[1030]);
  FullAdder FA1032 (Sum[933],Carry_out[977],Sum[978],Sum[1031],Carry_out[1031]);
  FullAdder FA1033 (Sum[934],Carry_out[978],Sum[979],Sum[1032],Carry_out[1032]);
  FullAdder FA1034 (Sum[935],Carry_out[979],Sum[980],Sum[1033],Carry_out[1033]);
  FullAdder FA1035 (Sum[936],Carry_out[980],Sum[981],Sum[1034],Carry_out[1034]);
  FullAdder FA1036 (Sum[937],Carry_out[981],Sum[982],Sum[1035],Carry_out[1035]);
  FullAdder FA1037 (Sum[938],Carry_out[982],Sum[983],Sum[1036],Carry_out[1036]);
  FullAdder FA1038 (Sum[939],Carry_out[983],Sum[984],Sum[1037],Carry_out[1037]);
  FullAdder FA1039 (Sum[940],Carry_out[984],Sum[985],Sum[1038],Carry_out[1038]);
  FullAdder FA1040 (Sum[941],Carry_out[985],Sum[986],Sum[1039],Carry_out[1039]);
  FullAdder FA1041 (Sum[942],Carry_out[986],Sum[987],Sum[1040],Carry_out[1040]);
  FullAdder FA1042 (Sum[943],Carry_out[987],Sum[988],Sum[1041],Carry_out[1041]);
  FullAdder FA1043 (Sum[944],Carry_out[988],Sum[989],Sum[1042],Carry_out[1042]);
  FullAdder FA1044 (Sum[945],Carry_out[989],Sum[990],Sum[1043],Carry_out[1043]);
  FullAdder FA1045 (Sum[946],Carry_out[990],Sum[991],Sum[1044],Carry_out[1044]);
  FullAdder FA1046 (Sum[947],Carry_out[991],Sum[992],Sum[1045],Carry_out[1045]);
  FullAdder FA1047 (Sum[948],Carry_out[992],Sum[993],Sum[1046],Carry_out[1046]);
  FullAdder FA1048 (Sum[949],Carry_out[993],Sum[994],Sum[1047],Carry_out[1047]);
  FullAdder FA1049 (Sum[950],Carry_out[994],Sum[995],Sum[1048],Carry_out[1048]);
  FullAdder FA1050 (Sum[951],Carry_out[995],Sum[996],Sum[1049],Carry_out[1049]);
  FullAdder FA1051 (Sum[952],Carry_out[996],Sum[997],Sum[1050],Carry_out[1050]);
  FullAdder FA1052 (Carry_out[952],Carry_out[997],Sum[998],Sum[1051],Carry_out[1051]);
  FullAdder FA1053 (Sum[900],Carry_out[998],Sum[999],Sum[1052],Carry_out[1052]);
  FullAdder FA1054 (Sum[901],Carry_out[999],Sum[1000],Sum[1053],Carry_out[1053]);
  FullAdder FA1055 (Sum[902],Carry_out[1000],Sum[1001],Sum[1054],Carry_out[1054]);
  FullAdder FA1056 (Sum[903],Carry_out[1001],Sum[1002],Sum[1055],Carry_out[1055]);
  FullAdder FA1057 (Sum[904],Carry_out[1002],Sum[1003],Sum[1056],Carry_out[1056]);
  FullAdder FA1058 (Sum[905],Carry_out[1003],Sum[1004],Sum[1057],Carry_out[1057]);
  FullAdder FA1059 (Sum[906],Carry_out[1004],Sum[1005],Sum[1058],Carry_out[1058]);
  FullAdder FA1060 (Carry_out[906],Carry_out[1005],Sum[1006],Sum[1059],Carry_out[1059]);
  FullAdder FA1061 (Carry_out[718],Sum[719],Carry_out[1006],Sum[1060],Carry_out[1060]);
  HalfAdder HA1062 (Partial_Product[31][31],Carry_out[719],Sum[1061],Carry_out[1061]);
  HalfAdder HA1063 (Carry_out[1007],Sum[1008],Sum[1062],Carry_out[1062]);
  FullAdder FA1064 (Carry_out[1008],Sum[1009],Carry_out[1062],Sum[1063],Carry_out[1063]);
  FullAdder FA1065 (Carry_out[1009],Sum[1010],Carry_out[1063],Sum[1064],Carry_out[1064]);
  FullAdder FA1066 (Carry_out[1010],Sum[1011],Carry_out[1064],Sum[1065],Carry_out[1065]);
  FullAdder FA1067 (Carry_out[1011],Sum[1012],Carry_out[1065],Sum[1066],Carry_out[1066]);
  FullAdder FA1068 (Carry_out[1012],Sum[1013],Carry_out[1066],Sum[1067],Carry_out[1067]);
  FullAdder FA1069 (Carry_out[1013],Sum[1014],Carry_out[1067],Sum[1068],Carry_out[1068]);
  FullAdder FA1070 (Carry_out[1014],Sum[1015],Carry_out[1068],Sum[1069],Carry_out[1069]);
  FullAdder FA1071 (Carry_out[1015],Sum[1016],Carry_out[1069],Sum[1070],Carry_out[1070]);
  FullAdder FA1072 (Carry_out[1016],Sum[1017],Carry_out[1070],Sum[1071],Carry_out[1071]);
  FullAdder FA1073 (Carry_out[1017],Sum[1018],Carry_out[1071],Sum[1072],Carry_out[1072]);
  FullAdder FA1074 (Carry_out[1018],Sum[1019],Carry_out[1072],Sum[1073],Carry_out[1073]);
  FullAdder FA1075 (Carry_out[1019],Sum[1020],Carry_out[1073],Sum[1074],Carry_out[1074]);
  FullAdder FA1076 (Carry_out[1020],Sum[1021],Carry_out[1074],Sum[1075],Carry_out[1075]);
  FullAdder FA1077 (Carry_out[1021],Sum[1022],Carry_out[1075],Sum[1076],Carry_out[1076]);
  FullAdder FA1078 (Carry_out[1022],Sum[1023],Carry_out[1076],Sum[1077],Carry_out[1077]);
  FullAdder FA1079 (Carry_out[1023],Sum[1024],Carry_out[1077],Sum[1078],Carry_out[1078]);
  FullAdder FA1080 (Carry_out[1024],Sum[1025],Carry_out[1078],Sum[1079],Carry_out[1079]);
  FullAdder FA1081 (Carry_out[1025],Sum[1026],Carry_out[1079],Sum[1080],Carry_out[1080]);
  FullAdder FA1082 (Carry_out[1026],Sum[1027],Carry_out[1080],Sum[1081],Carry_out[1081]);
  FullAdder FA1083 (Carry_out[1027],Sum[1028],Carry_out[1081],Sum[1082],Carry_out[1082]);
  FullAdder FA1084 (Carry_out[1028],Sum[1029],Carry_out[1082],Sum[1083],Carry_out[1083]);
  FullAdder FA1085 (Carry_out[1029],Sum[1030],Carry_out[1083],Sum[1084],Carry_out[1084]);
  FullAdder FA1086 (Carry_out[1030],Sum[1031],Carry_out[1084],Sum[1085],Carry_out[1085]);
  FullAdder FA1087 (Carry_out[1031],Sum[1032],Carry_out[1085],Sum[1086],Carry_out[1086]);
  FullAdder FA1088 (Carry_out[1032],Sum[1033],Carry_out[1086],Sum[1087],Carry_out[1087]);
  FullAdder FA1089 (Carry_out[1033],Sum[1034],Carry_out[1087],Sum[1088],Carry_out[1088]);
  FullAdder FA1090 (Carry_out[1034],Sum[1035],Carry_out[1088],Sum[1089],Carry_out[1089]);
  FullAdder FA1091 (Carry_out[1035],Sum[1036],Carry_out[1089],Sum[1090],Carry_out[1090]);
  FullAdder FA1092 (Carry_out[1036],Sum[1037],Carry_out[1090],Sum[1091],Carry_out[1091]);
  FullAdder FA1093 (Carry_out[1037],Sum[1038],Carry_out[1091],Sum[1092],Carry_out[1092]);
  FullAdder FA1094 (Carry_out[1038],Sum[1039],Carry_out[1092],Sum[1093],Carry_out[1093]);
  FullAdder FA1095 (Carry_out[1039],Sum[1040],Carry_out[1093],Sum[1094],Carry_out[1094]);
  FullAdder FA1096 (Carry_out[1040],Sum[1041],Carry_out[1094],Sum[1095],Carry_out[1095]);
  FullAdder FA1097 (Carry_out[1041],Sum[1042],Carry_out[1095],Sum[1096],Carry_out[1096]);
  FullAdder FA1098 (Carry_out[1042],Sum[1043],Carry_out[1096],Sum[1097],Carry_out[1097]);
  FullAdder FA1099 (Carry_out[1043],Sum[1044],Carry_out[1097],Sum[1098],Carry_out[1098]);
  FullAdder FA1100 (Carry_out[1044],Sum[1045],Carry_out[1098],Sum[1099],Carry_out[1099]);
  FullAdder FA1101 (Carry_out[1045],Sum[1046],Carry_out[1099],Sum[1100],Carry_out[1100]);
  FullAdder FA1102 (Carry_out[1046],Sum[1047],Carry_out[1100],Sum[1101],Carry_out[1101]);
  FullAdder FA1103 (Carry_out[1047],Sum[1048],Carry_out[1101],Sum[1102],Carry_out[1102]);
  FullAdder FA1104 (Carry_out[1048],Sum[1049],Carry_out[1102],Sum[1103],Carry_out[1103]);
  FullAdder FA1105 (Carry_out[1049],Sum[1050],Carry_out[1103],Sum[1104],Carry_out[1104]);
  FullAdder FA1106 (Carry_out[1050],Sum[1051],Carry_out[1104],Sum[1105],Carry_out[1105]);
  FullAdder FA1107 (Carry_out[1051],Sum[1052],Carry_out[1105],Sum[1106],Carry_out[1106]);
  FullAdder FA1108 (Carry_out[1052],Sum[1053],Carry_out[1106],Sum[1107],Carry_out[1107]);
  FullAdder FA1109 (Carry_out[1053],Sum[1054],Carry_out[1107],Sum[1108],Carry_out[1108]);
  FullAdder FA1110 (Carry_out[1054],Sum[1055],Carry_out[1108],Sum[1109],Carry_out[1109]);
  FullAdder FA1111 (Carry_out[1055],Sum[1056],Carry_out[1109],Sum[1110],Carry_out[1110]);
  FullAdder FA1112 (Carry_out[1056],Sum[1057],Carry_out[1110],Sum[1111],Carry_out[1111]);
  FullAdder FA1113 (Carry_out[1057],Sum[1058],Carry_out[1111],Sum[1112],Carry_out[1112]);
  FullAdder FA1114 (Carry_out[1058],Sum[1059],Carry_out[1112],Sum[1113],Carry_out[1113]);
  FullAdder FA1115 (Carry_out[1059],Sum[1060],Carry_out[1113],Sum[1114],Carry_out[1114]);
  FullAdder FA1116 (Carry_out[1060],Sum[1061],Carry_out[1114],Sum[1115],Carry_out[1115]);
  HalfAdder HA1117 (Carry_out[1061],Carry_out[1115],Sum[1116],Carry_out[1116]);



//Assigning final Sum to the Final product bit wise
//we can also use concatination operator
  assign Final_Product[63] = Sum[1116];
  assign Final_Product[62] = Sum[1115];
  assign Final_Product[61] = Sum[1114];
  assign Final_Product[60] = Sum[1113];
  assign Final_Product[59] = Sum[1112];
  assign Final_Product[58] = Sum[1111];
  assign Final_Product[57] = Sum[1110];
  assign Final_Product[56] = Sum[1109];
  assign Final_Product[55] = Sum[1108];
  assign Final_Product[54] = Sum[1107];
  assign Final_Product[53] = Sum[1106];
  assign Final_Product[52] = Sum[1105];
  assign Final_Product[51] = Sum[1104];
  assign Final_Product[50] = Sum[1103];
  assign Final_Product[49] = Sum[1102];
  assign Final_Product[48] = Sum[1101];
  assign Final_Product[47] = Sum[1100];
  assign Final_Product[46] = Sum[1099];
  assign Final_Product[45] = Sum[1098];
  assign Final_Product[44] = Sum[1097];
  assign Final_Product[43] = Sum[1096];
  assign Final_Product[42] = Sum[1095];
  assign Final_Product[41] = Sum[1094];
  assign Final_Product[40] = Sum[1093];
  assign Final_Product[39] = Sum[1092];
  assign Final_Product[38] = Sum[1091];
  assign Final_Product[37] = Sum[1090];
  assign Final_Product[36] = Sum[1089];
  assign Final_Product[35] = Sum[1088];
  assign Final_Product[34] = Sum[1087];
  assign Final_Product[33] = Sum[1086];
  assign Final_Product[32] = Sum[1085];
  assign Final_Product[31] = Sum[1084];
  assign Final_Product[30] = Sum[1083];
  assign Final_Product[29] = Sum[1082];
  assign Final_Product[28] = Sum[1081];
  assign Final_Product[27] = Sum[1080];
  assign Final_Product[26] = Sum[1079];
  assign Final_Product[25] = Sum[1078];
  assign Final_Product[24] = Sum[1077];
  assign Final_Product[23] = Sum[1076];
  assign Final_Product[22] = Sum[1075];
  assign Final_Product[21] = Sum[1074];
  assign Final_Product[20] = Sum[1073];
  assign Final_Product[19] = Sum[1072];
  assign Final_Product[18] = Sum[1071];
  assign Final_Product[17] = Sum[1070];
  assign Final_Product[16] = Sum[1069];
  assign Final_Product[15] = Sum[1068];
  assign Final_Product[14] = Sum[1067];
  assign Final_Product[13] = Sum[1066];
  assign Final_Product[12] = Sum[1065];
  assign Final_Product[11] = Sum[1064];
  assign Final_Product[10] = Sum[1063];
  assign Final_Product[9]  = Sum[1062];
  assign Final_Product[8]  = Sum[1007];
  assign Final_Product[7]  = Sum[953];
  assign Final_Product[6]  = Sum[907];
  assign Final_Product[5]  = Sum[828];
  assign Final_Product[4]  = Sum[720];
  assign Final_Product[3]  = Sum[550];
  assign Final_Product[2]  = Sum[320];
  assign Final_Product[1]  = Sum[0];
  assign Final_Product[0]  = Partial_Product[0][0];
endmodule

