`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2024 Talha Mahboob
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
///////////////////////////////////////////////////////////////////////////////

module ModularReduction (
  input  logic [255:0] in ,
  output logic [127:0] out
);

  // Polynomial for GF(2^128)
  localparam logic [127:0] POLY = 128'hE1000000000000000000000000000000;

  logic [255:0] temp;
  logic [127:0] high, low;

  // Initial assignment
  assign temp = in;

  // Reduction process
  always_comb begin
    high = temp[255:128];
    low  = temp[127:0];

    // Perform reduction
    for (int i = 127; i >= 0; i--) begin
      if (high[i]) begin
        high = high ^ (POLY << (i - 128));
        low  = low ^ (POLY << (i - 128));
      end
    end

    out = low;
  end
endmodule